module InstFetch(
  input         clock,
  input         reset,
  output        io_imem_inst_valid,
  input         io_imem_inst_ready,
  output [31:0] io_imem_inst_addr,
  input  [31:0] io_imem_inst_read,
  input  [1:0]  io_pcSrc,
  input  [31:0] io_nextPC,
  input         io_stall,
  input         io_memDone,
  output        io_out_valid,
  output [31:0] io_out_pc,
  output [31:0] io_out_inst,
  output        io_IFDone
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] pc; // @[InstFetch.scala 29:19]
  reg [31:0] inst; // @[InstFetch.scala 30:21]
  wire  _io_imem_inst_valid_T = ~io_stall; // @[InstFetch.scala 32:25]
  wire  _fire_T = io_imem_inst_valid & io_imem_inst_ready; // @[InstFetch.scala 38:34]
  wire  fire = io_stall | _fire_T; // @[InstFetch.scala 37:17]
  reg  ifPCfire; // @[InstFetch.scala 41:25]
  reg  ifPCstall; // @[InstFetch.scala 42:26]
  wire [31:0] _ifPC_T_4 = pc + 32'h4; // @[InstFetch.scala 44:40]
  wire [31:0] _ifPC_T_5 = io_pcSrc == 2'h0 ? _ifPC_T_4 : io_nextPC; // @[InstFetch.scala 44:18]
  assign io_imem_inst_valid = ~io_stall; // @[InstFetch.scala 32:25]
  assign io_imem_inst_addr = pc; // @[InstFetch.scala 34:21]
  assign io_out_valid = io_stall | _fire_T; // @[InstFetch.scala 37:17]
  assign io_out_pc = ifPCfire & ~ifPCstall ? _ifPC_T_5 : pc; // @[InstFetch.scala 43:17]
  assign io_out_inst = fire & _io_imem_inst_valid_T ? io_imem_inst_read : inst; // @[InstFetch.scala 40:19]
  assign io_IFDone = fire & io_memDone; // @[InstFetch.scala 50:21]
  always @(posedge clock) begin
    if (reset) begin // @[InstFetch.scala 29:19]
      pc <= 32'h80000000; // @[InstFetch.scala 29:19]
    end else if (ifPCfire & ~ifPCstall) begin // @[InstFetch.scala 43:17]
      if (io_pcSrc == 2'h0) begin // @[InstFetch.scala 44:18]
        pc <= _ifPC_T_4;
      end else begin
        pc <= io_nextPC;
      end
    end
    if (reset) begin // @[InstFetch.scala 30:21]
      inst <= 32'h0; // @[InstFetch.scala 30:21]
    end else if (fire & _io_imem_inst_valid_T) begin // @[InstFetch.scala 40:19]
      inst <= io_imem_inst_read;
    end
    ifPCfire <= io_stall | _fire_T; // @[InstFetch.scala 37:17]
    ifPCstall <= io_stall; // @[InstFetch.scala 42:26]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  pc = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  inst = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  ifPCfire = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  ifPCstall = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PipelineReg(
  input         clock,
  input         reset,
  input         io_in_valid,
  input  [31:0] io_in_pc,
  input  [31:0] io_in_inst,
  input         io_in_typeL,
  input         io_in_aluA,
  input  [1:0]  io_in_aluB,
  input  [3:0]  io_in_aluOp,
  input  [2:0]  io_in_branch,
  input  [1:0]  io_in_memtoReg,
  input         io_in_memWr,
  input  [2:0]  io_in_memOp,
  input         io_in_rdEn,
  input  [4:0]  io_in_rdAddr,
  input  [63:0] io_in_rs1Data,
  input  [63:0] io_in_rs2Data,
  input  [63:0] io_in_imm,
  input  [63:0] io_in_aluRes,
  input  [63:0] io_in_memData,
  output        io_out_valid,
  output [31:0] io_out_pc,
  output [31:0] io_out_inst,
  output        io_out_typeL,
  output        io_out_aluA,
  output [1:0]  io_out_aluB,
  output [3:0]  io_out_aluOp,
  output [2:0]  io_out_branch,
  output [1:0]  io_out_memtoReg,
  output        io_out_memWr,
  output [2:0]  io_out_memOp,
  output        io_out_rdEn,
  output [4:0]  io_out_rdAddr,
  output [63:0] io_out_rs1Data,
  output [63:0] io_out_rs2Data,
  output [63:0] io_out_imm,
  output [63:0] io_out_aluRes,
  output [63:0] io_out_memData,
  input         io_flush,
  input         io_stall
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
`endif // RANDOMIZE_REG_INIT
  reg  reg_valid; // @[PipelineReg.scala 75:20]
  reg [31:0] reg_pc; // @[PipelineReg.scala 75:20]
  reg [31:0] reg_inst; // @[PipelineReg.scala 75:20]
  reg  reg_typeL; // @[PipelineReg.scala 75:20]
  reg  reg_aluA; // @[PipelineReg.scala 75:20]
  reg [1:0] reg_aluB; // @[PipelineReg.scala 75:20]
  reg [3:0] reg_aluOp; // @[PipelineReg.scala 75:20]
  reg [2:0] reg_branch; // @[PipelineReg.scala 75:20]
  reg [1:0] reg_memtoReg; // @[PipelineReg.scala 75:20]
  reg  reg_memWr; // @[PipelineReg.scala 75:20]
  reg [2:0] reg_memOp; // @[PipelineReg.scala 75:20]
  reg  reg_rdEn; // @[PipelineReg.scala 75:20]
  reg [4:0] reg_rdAddr; // @[PipelineReg.scala 75:20]
  reg [63:0] reg_rs1Data; // @[PipelineReg.scala 75:20]
  reg [63:0] reg_rs2Data; // @[PipelineReg.scala 75:20]
  reg [63:0] reg_imm; // @[PipelineReg.scala 75:20]
  reg [63:0] reg_aluRes; // @[PipelineReg.scala 75:20]
  reg [63:0] reg_memData; // @[PipelineReg.scala 75:20]
  wire  _T = ~io_stall; // @[PipelineReg.scala 77:33]
  assign io_out_valid = reg_valid; // @[PipelineReg.scala 83:10]
  assign io_out_pc = reg_pc; // @[PipelineReg.scala 83:10]
  assign io_out_inst = reg_inst; // @[PipelineReg.scala 83:10]
  assign io_out_typeL = reg_typeL; // @[PipelineReg.scala 83:10]
  assign io_out_aluA = reg_aluA; // @[PipelineReg.scala 83:10]
  assign io_out_aluB = reg_aluB; // @[PipelineReg.scala 83:10]
  assign io_out_aluOp = reg_aluOp; // @[PipelineReg.scala 83:10]
  assign io_out_branch = reg_branch; // @[PipelineReg.scala 83:10]
  assign io_out_memtoReg = reg_memtoReg; // @[PipelineReg.scala 83:10]
  assign io_out_memWr = reg_memWr; // @[PipelineReg.scala 83:10]
  assign io_out_memOp = reg_memOp; // @[PipelineReg.scala 83:10]
  assign io_out_rdEn = reg_rdEn; // @[PipelineReg.scala 83:10]
  assign io_out_rdAddr = reg_rdAddr; // @[PipelineReg.scala 83:10]
  assign io_out_rs1Data = reg_rs1Data; // @[PipelineReg.scala 83:10]
  assign io_out_rs2Data = reg_rs2Data; // @[PipelineReg.scala 83:10]
  assign io_out_imm = reg_imm; // @[PipelineReg.scala 83:10]
  assign io_out_aluRes = reg_aluRes; // @[PipelineReg.scala 83:10]
  assign io_out_memData = reg_memData; // @[PipelineReg.scala 83:10]
  always @(posedge clock) begin
    if (reset) begin // @[PipelineReg.scala 75:20]
      reg_valid <= 1'h0; // @[PipelineReg.scala 75:20]
    end else if (io_flush & ~io_stall) begin // @[PipelineReg.scala 77:44]
      reg_valid <= 1'h0; // @[PipelineReg.scala 34:14]
    end else if (_T) begin // @[PipelineReg.scala 79:27]
      reg_valid <= io_in_valid; // @[PipelineReg.scala 80:9]
    end
    if (reset) begin // @[PipelineReg.scala 75:20]
      reg_pc <= 32'h0; // @[PipelineReg.scala 75:20]
    end else if (io_flush & ~io_stall) begin // @[PipelineReg.scala 77:44]
      reg_pc <= 32'h0; // @[PipelineReg.scala 35:14]
    end else if (_T) begin // @[PipelineReg.scala 79:27]
      reg_pc <= io_in_pc; // @[PipelineReg.scala 80:9]
    end
    if (reset) begin // @[PipelineReg.scala 75:20]
      reg_inst <= 32'h0; // @[PipelineReg.scala 75:20]
    end else if (io_flush & ~io_stall) begin // @[PipelineReg.scala 77:44]
      reg_inst <= 32'h0; // @[PipelineReg.scala 36:14]
    end else if (_T) begin // @[PipelineReg.scala 79:27]
      reg_inst <= io_in_inst; // @[PipelineReg.scala 80:9]
    end
    if (reset) begin // @[PipelineReg.scala 75:20]
      reg_typeL <= 1'h0; // @[PipelineReg.scala 75:20]
    end else if (io_flush & ~io_stall) begin // @[PipelineReg.scala 77:44]
      reg_typeL <= 1'h0; // @[PipelineReg.scala 37:14]
    end else if (_T) begin // @[PipelineReg.scala 79:27]
      reg_typeL <= io_in_typeL; // @[PipelineReg.scala 80:9]
    end
    if (reset) begin // @[PipelineReg.scala 75:20]
      reg_aluA <= 1'h0; // @[PipelineReg.scala 75:20]
    end else if (io_flush & ~io_stall) begin // @[PipelineReg.scala 77:44]
      reg_aluA <= 1'h0; // @[PipelineReg.scala 39:14]
    end else if (_T) begin // @[PipelineReg.scala 79:27]
      reg_aluA <= io_in_aluA; // @[PipelineReg.scala 80:9]
    end
    if (reset) begin // @[PipelineReg.scala 75:20]
      reg_aluB <= 2'h0; // @[PipelineReg.scala 75:20]
    end else if (io_flush & ~io_stall) begin // @[PipelineReg.scala 77:44]
      reg_aluB <= 2'h3; // @[PipelineReg.scala 40:14]
    end else if (_T) begin // @[PipelineReg.scala 79:27]
      reg_aluB <= io_in_aluB; // @[PipelineReg.scala 80:9]
    end
    if (reset) begin // @[PipelineReg.scala 75:20]
      reg_aluOp <= 4'h0; // @[PipelineReg.scala 75:20]
    end else if (io_flush & ~io_stall) begin // @[PipelineReg.scala 77:44]
      reg_aluOp <= 4'h0; // @[PipelineReg.scala 41:14]
    end else if (_T) begin // @[PipelineReg.scala 79:27]
      reg_aluOp <= io_in_aluOp; // @[PipelineReg.scala 80:9]
    end
    if (reset) begin // @[PipelineReg.scala 75:20]
      reg_branch <= 3'h0; // @[PipelineReg.scala 75:20]
    end else if (io_flush & ~io_stall) begin // @[PipelineReg.scala 77:44]
      reg_branch <= 3'h0; // @[PipelineReg.scala 43:14]
    end else if (_T) begin // @[PipelineReg.scala 79:27]
      reg_branch <= io_in_branch; // @[PipelineReg.scala 80:9]
    end
    if (reset) begin // @[PipelineReg.scala 75:20]
      reg_memtoReg <= 2'h0; // @[PipelineReg.scala 75:20]
    end else if (io_flush & ~io_stall) begin // @[PipelineReg.scala 77:44]
      reg_memtoReg <= 2'h0; // @[PipelineReg.scala 44:14]
    end else if (_T) begin // @[PipelineReg.scala 79:27]
      reg_memtoReg <= io_in_memtoReg; // @[PipelineReg.scala 80:9]
    end
    if (reset) begin // @[PipelineReg.scala 75:20]
      reg_memWr <= 1'h0; // @[PipelineReg.scala 75:20]
    end else if (io_flush & ~io_stall) begin // @[PipelineReg.scala 77:44]
      reg_memWr <= 1'h0; // @[PipelineReg.scala 45:14]
    end else if (_T) begin // @[PipelineReg.scala 79:27]
      reg_memWr <= io_in_memWr; // @[PipelineReg.scala 80:9]
    end
    if (reset) begin // @[PipelineReg.scala 75:20]
      reg_memOp <= 3'h0; // @[PipelineReg.scala 75:20]
    end else if (io_flush & ~io_stall) begin // @[PipelineReg.scala 77:44]
      reg_memOp <= 3'h0; // @[PipelineReg.scala 46:14]
    end else if (_T) begin // @[PipelineReg.scala 79:27]
      reg_memOp <= io_in_memOp; // @[PipelineReg.scala 80:9]
    end
    if (reset) begin // @[PipelineReg.scala 75:20]
      reg_rdEn <= 1'h0; // @[PipelineReg.scala 75:20]
    end else if (io_flush & ~io_stall) begin // @[PipelineReg.scala 77:44]
      reg_rdEn <= 1'h0; // @[PipelineReg.scala 48:14]
    end else if (_T) begin // @[PipelineReg.scala 79:27]
      reg_rdEn <= io_in_rdEn; // @[PipelineReg.scala 80:9]
    end
    if (reset) begin // @[PipelineReg.scala 75:20]
      reg_rdAddr <= 5'h0; // @[PipelineReg.scala 75:20]
    end else if (io_flush & ~io_stall) begin // @[PipelineReg.scala 77:44]
      reg_rdAddr <= 5'h0; // @[PipelineReg.scala 49:14]
    end else if (_T) begin // @[PipelineReg.scala 79:27]
      reg_rdAddr <= io_in_rdAddr; // @[PipelineReg.scala 80:9]
    end
    if (reset) begin // @[PipelineReg.scala 75:20]
      reg_rs1Data <= 64'h0; // @[PipelineReg.scala 75:20]
    end else if (io_flush & ~io_stall) begin // @[PipelineReg.scala 77:44]
      reg_rs1Data <= 64'h0; // @[PipelineReg.scala 51:14]
    end else if (_T) begin // @[PipelineReg.scala 79:27]
      reg_rs1Data <= io_in_rs1Data; // @[PipelineReg.scala 80:9]
    end
    if (reset) begin // @[PipelineReg.scala 75:20]
      reg_rs2Data <= 64'h0; // @[PipelineReg.scala 75:20]
    end else if (io_flush & ~io_stall) begin // @[PipelineReg.scala 77:44]
      reg_rs2Data <= 64'h0; // @[PipelineReg.scala 52:14]
    end else if (_T) begin // @[PipelineReg.scala 79:27]
      reg_rs2Data <= io_in_rs2Data; // @[PipelineReg.scala 80:9]
    end
    if (reset) begin // @[PipelineReg.scala 75:20]
      reg_imm <= 64'h0; // @[PipelineReg.scala 75:20]
    end else if (io_flush & ~io_stall) begin // @[PipelineReg.scala 77:44]
      reg_imm <= 64'h0; // @[PipelineReg.scala 53:14]
    end else if (_T) begin // @[PipelineReg.scala 79:27]
      reg_imm <= io_in_imm; // @[PipelineReg.scala 80:9]
    end
    if (reset) begin // @[PipelineReg.scala 75:20]
      reg_aluRes <= 64'h0; // @[PipelineReg.scala 75:20]
    end else if (io_flush & ~io_stall) begin // @[PipelineReg.scala 77:44]
      reg_aluRes <= 64'h0; // @[PipelineReg.scala 57:14]
    end else if (_T) begin // @[PipelineReg.scala 79:27]
      reg_aluRes <= io_in_aluRes; // @[PipelineReg.scala 80:9]
    end
    if (reset) begin // @[PipelineReg.scala 75:20]
      reg_memData <= 64'h0; // @[PipelineReg.scala 75:20]
    end else if (io_flush & ~io_stall) begin // @[PipelineReg.scala 77:44]
      reg_memData <= 64'h0; // @[PipelineReg.scala 58:16]
    end else if (_T) begin // @[PipelineReg.scala 79:27]
      reg_memData <= io_in_memData; // @[PipelineReg.scala 80:9]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reg_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  reg_pc = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  reg_inst = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  reg_typeL = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  reg_aluA = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  reg_aluB = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  reg_aluOp = _RAND_6[3:0];
  _RAND_7 = {1{`RANDOM}};
  reg_branch = _RAND_7[2:0];
  _RAND_8 = {1{`RANDOM}};
  reg_memtoReg = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  reg_memWr = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  reg_memOp = _RAND_10[2:0];
  _RAND_11 = {1{`RANDOM}};
  reg_rdEn = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  reg_rdAddr = _RAND_12[4:0];
  _RAND_13 = {2{`RANDOM}};
  reg_rs1Data = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  reg_rs2Data = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  reg_imm = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  reg_aluRes = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  reg_memData = _RAND_17[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RegFile(
  input         clock,
  input         reset,
  output [63:0] io_rs1Data,
  output [63:0] io_rs2Data,
  input         io_rdEn,
  input  [31:0] io_rdAddr,
  input  [63:0] io_rdData,
  input         io_ctrl_rs1En,
  input         io_ctrl_rs2En,
  input  [4:0]  io_ctrl_rs1Addr,
  input  [4:0]  io_ctrl_rs2Addr,
  output [63:0] rf_10
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
`endif // RANDOMIZE_REG_INIT
  wire  dt_ar_clock; // @[RegFile.scala 26:21]
  wire [7:0] dt_ar_coreid; // @[RegFile.scala 26:21]
  wire [63:0] dt_ar_gpr_0; // @[RegFile.scala 26:21]
  wire [63:0] dt_ar_gpr_1; // @[RegFile.scala 26:21]
  wire [63:0] dt_ar_gpr_2; // @[RegFile.scala 26:21]
  wire [63:0] dt_ar_gpr_3; // @[RegFile.scala 26:21]
  wire [63:0] dt_ar_gpr_4; // @[RegFile.scala 26:21]
  wire [63:0] dt_ar_gpr_5; // @[RegFile.scala 26:21]
  wire [63:0] dt_ar_gpr_6; // @[RegFile.scala 26:21]
  wire [63:0] dt_ar_gpr_7; // @[RegFile.scala 26:21]
  wire [63:0] dt_ar_gpr_8; // @[RegFile.scala 26:21]
  wire [63:0] dt_ar_gpr_9; // @[RegFile.scala 26:21]
  wire [63:0] dt_ar_gpr_10; // @[RegFile.scala 26:21]
  wire [63:0] dt_ar_gpr_11; // @[RegFile.scala 26:21]
  wire [63:0] dt_ar_gpr_12; // @[RegFile.scala 26:21]
  wire [63:0] dt_ar_gpr_13; // @[RegFile.scala 26:21]
  wire [63:0] dt_ar_gpr_14; // @[RegFile.scala 26:21]
  wire [63:0] dt_ar_gpr_15; // @[RegFile.scala 26:21]
  wire [63:0] dt_ar_gpr_16; // @[RegFile.scala 26:21]
  wire [63:0] dt_ar_gpr_17; // @[RegFile.scala 26:21]
  wire [63:0] dt_ar_gpr_18; // @[RegFile.scala 26:21]
  wire [63:0] dt_ar_gpr_19; // @[RegFile.scala 26:21]
  wire [63:0] dt_ar_gpr_20; // @[RegFile.scala 26:21]
  wire [63:0] dt_ar_gpr_21; // @[RegFile.scala 26:21]
  wire [63:0] dt_ar_gpr_22; // @[RegFile.scala 26:21]
  wire [63:0] dt_ar_gpr_23; // @[RegFile.scala 26:21]
  wire [63:0] dt_ar_gpr_24; // @[RegFile.scala 26:21]
  wire [63:0] dt_ar_gpr_25; // @[RegFile.scala 26:21]
  wire [63:0] dt_ar_gpr_26; // @[RegFile.scala 26:21]
  wire [63:0] dt_ar_gpr_27; // @[RegFile.scala 26:21]
  wire [63:0] dt_ar_gpr_28; // @[RegFile.scala 26:21]
  wire [63:0] dt_ar_gpr_29; // @[RegFile.scala 26:21]
  wire [63:0] dt_ar_gpr_30; // @[RegFile.scala 26:21]
  wire [63:0] dt_ar_gpr_31; // @[RegFile.scala 26:21]
  reg [63:0] rf__0; // @[RegFile.scala 17:19]
  reg [63:0] rf__1; // @[RegFile.scala 17:19]
  reg [63:0] rf__2; // @[RegFile.scala 17:19]
  reg [63:0] rf__3; // @[RegFile.scala 17:19]
  reg [63:0] rf__4; // @[RegFile.scala 17:19]
  reg [63:0] rf__5; // @[RegFile.scala 17:19]
  reg [63:0] rf__6; // @[RegFile.scala 17:19]
  reg [63:0] rf__7; // @[RegFile.scala 17:19]
  reg [63:0] rf__8; // @[RegFile.scala 17:19]
  reg [63:0] rf__9; // @[RegFile.scala 17:19]
  reg [63:0] rf__10; // @[RegFile.scala 17:19]
  reg [63:0] rf__11; // @[RegFile.scala 17:19]
  reg [63:0] rf__12; // @[RegFile.scala 17:19]
  reg [63:0] rf__13; // @[RegFile.scala 17:19]
  reg [63:0] rf__14; // @[RegFile.scala 17:19]
  reg [63:0] rf__15; // @[RegFile.scala 17:19]
  reg [63:0] rf__16; // @[RegFile.scala 17:19]
  reg [63:0] rf__17; // @[RegFile.scala 17:19]
  reg [63:0] rf__18; // @[RegFile.scala 17:19]
  reg [63:0] rf__19; // @[RegFile.scala 17:19]
  reg [63:0] rf__20; // @[RegFile.scala 17:19]
  reg [63:0] rf__21; // @[RegFile.scala 17:19]
  reg [63:0] rf__22; // @[RegFile.scala 17:19]
  reg [63:0] rf__23; // @[RegFile.scala 17:19]
  reg [63:0] rf__24; // @[RegFile.scala 17:19]
  reg [63:0] rf__25; // @[RegFile.scala 17:19]
  reg [63:0] rf__26; // @[RegFile.scala 17:19]
  reg [63:0] rf__27; // @[RegFile.scala 17:19]
  reg [63:0] rf__28; // @[RegFile.scala 17:19]
  reg [63:0] rf__29; // @[RegFile.scala 17:19]
  reg [63:0] rf__30; // @[RegFile.scala 17:19]
  reg [63:0] rf__31; // @[RegFile.scala 17:19]
  wire [63:0] _GEN_65 = 5'h1 == io_ctrl_rs1Addr ? rf__1 : rf__0; // @[RegFile.scala 23:{20,20}]
  wire [63:0] _GEN_66 = 5'h2 == io_ctrl_rs1Addr ? rf__2 : _GEN_65; // @[RegFile.scala 23:{20,20}]
  wire [63:0] _GEN_67 = 5'h3 == io_ctrl_rs1Addr ? rf__3 : _GEN_66; // @[RegFile.scala 23:{20,20}]
  wire [63:0] _GEN_68 = 5'h4 == io_ctrl_rs1Addr ? rf__4 : _GEN_67; // @[RegFile.scala 23:{20,20}]
  wire [63:0] _GEN_69 = 5'h5 == io_ctrl_rs1Addr ? rf__5 : _GEN_68; // @[RegFile.scala 23:{20,20}]
  wire [63:0] _GEN_70 = 5'h6 == io_ctrl_rs1Addr ? rf__6 : _GEN_69; // @[RegFile.scala 23:{20,20}]
  wire [63:0] _GEN_71 = 5'h7 == io_ctrl_rs1Addr ? rf__7 : _GEN_70; // @[RegFile.scala 23:{20,20}]
  wire [63:0] _GEN_72 = 5'h8 == io_ctrl_rs1Addr ? rf__8 : _GEN_71; // @[RegFile.scala 23:{20,20}]
  wire [63:0] _GEN_73 = 5'h9 == io_ctrl_rs1Addr ? rf__9 : _GEN_72; // @[RegFile.scala 23:{20,20}]
  wire [63:0] _GEN_74 = 5'ha == io_ctrl_rs1Addr ? rf__10 : _GEN_73; // @[RegFile.scala 23:{20,20}]
  wire [63:0] _GEN_75 = 5'hb == io_ctrl_rs1Addr ? rf__11 : _GEN_74; // @[RegFile.scala 23:{20,20}]
  wire [63:0] _GEN_76 = 5'hc == io_ctrl_rs1Addr ? rf__12 : _GEN_75; // @[RegFile.scala 23:{20,20}]
  wire [63:0] _GEN_77 = 5'hd == io_ctrl_rs1Addr ? rf__13 : _GEN_76; // @[RegFile.scala 23:{20,20}]
  wire [63:0] _GEN_78 = 5'he == io_ctrl_rs1Addr ? rf__14 : _GEN_77; // @[RegFile.scala 23:{20,20}]
  wire [63:0] _GEN_79 = 5'hf == io_ctrl_rs1Addr ? rf__15 : _GEN_78; // @[RegFile.scala 23:{20,20}]
  wire [63:0] _GEN_80 = 5'h10 == io_ctrl_rs1Addr ? rf__16 : _GEN_79; // @[RegFile.scala 23:{20,20}]
  wire [63:0] _GEN_81 = 5'h11 == io_ctrl_rs1Addr ? rf__17 : _GEN_80; // @[RegFile.scala 23:{20,20}]
  wire [63:0] _GEN_82 = 5'h12 == io_ctrl_rs1Addr ? rf__18 : _GEN_81; // @[RegFile.scala 23:{20,20}]
  wire [63:0] _GEN_83 = 5'h13 == io_ctrl_rs1Addr ? rf__19 : _GEN_82; // @[RegFile.scala 23:{20,20}]
  wire [63:0] _GEN_84 = 5'h14 == io_ctrl_rs1Addr ? rf__20 : _GEN_83; // @[RegFile.scala 23:{20,20}]
  wire [63:0] _GEN_85 = 5'h15 == io_ctrl_rs1Addr ? rf__21 : _GEN_84; // @[RegFile.scala 23:{20,20}]
  wire [63:0] _GEN_86 = 5'h16 == io_ctrl_rs1Addr ? rf__22 : _GEN_85; // @[RegFile.scala 23:{20,20}]
  wire [63:0] _GEN_87 = 5'h17 == io_ctrl_rs1Addr ? rf__23 : _GEN_86; // @[RegFile.scala 23:{20,20}]
  wire [63:0] _GEN_88 = 5'h18 == io_ctrl_rs1Addr ? rf__24 : _GEN_87; // @[RegFile.scala 23:{20,20}]
  wire [63:0] _GEN_89 = 5'h19 == io_ctrl_rs1Addr ? rf__25 : _GEN_88; // @[RegFile.scala 23:{20,20}]
  wire [63:0] _GEN_90 = 5'h1a == io_ctrl_rs1Addr ? rf__26 : _GEN_89; // @[RegFile.scala 23:{20,20}]
  wire [63:0] _GEN_91 = 5'h1b == io_ctrl_rs1Addr ? rf__27 : _GEN_90; // @[RegFile.scala 23:{20,20}]
  wire [63:0] _GEN_92 = 5'h1c == io_ctrl_rs1Addr ? rf__28 : _GEN_91; // @[RegFile.scala 23:{20,20}]
  wire [63:0] _GEN_93 = 5'h1d == io_ctrl_rs1Addr ? rf__29 : _GEN_92; // @[RegFile.scala 23:{20,20}]
  wire [63:0] _GEN_94 = 5'h1e == io_ctrl_rs1Addr ? rf__30 : _GEN_93; // @[RegFile.scala 23:{20,20}]
  wire [63:0] _GEN_95 = 5'h1f == io_ctrl_rs1Addr ? rf__31 : _GEN_94; // @[RegFile.scala 23:{20,20}]
  wire [63:0] _GEN_97 = 5'h1 == io_ctrl_rs2Addr ? rf__1 : rf__0; // @[RegFile.scala 24:{20,20}]
  wire [63:0] _GEN_98 = 5'h2 == io_ctrl_rs2Addr ? rf__2 : _GEN_97; // @[RegFile.scala 24:{20,20}]
  wire [63:0] _GEN_99 = 5'h3 == io_ctrl_rs2Addr ? rf__3 : _GEN_98; // @[RegFile.scala 24:{20,20}]
  wire [63:0] _GEN_100 = 5'h4 == io_ctrl_rs2Addr ? rf__4 : _GEN_99; // @[RegFile.scala 24:{20,20}]
  wire [63:0] _GEN_101 = 5'h5 == io_ctrl_rs2Addr ? rf__5 : _GEN_100; // @[RegFile.scala 24:{20,20}]
  wire [63:0] _GEN_102 = 5'h6 == io_ctrl_rs2Addr ? rf__6 : _GEN_101; // @[RegFile.scala 24:{20,20}]
  wire [63:0] _GEN_103 = 5'h7 == io_ctrl_rs2Addr ? rf__7 : _GEN_102; // @[RegFile.scala 24:{20,20}]
  wire [63:0] _GEN_104 = 5'h8 == io_ctrl_rs2Addr ? rf__8 : _GEN_103; // @[RegFile.scala 24:{20,20}]
  wire [63:0] _GEN_105 = 5'h9 == io_ctrl_rs2Addr ? rf__9 : _GEN_104; // @[RegFile.scala 24:{20,20}]
  wire [63:0] _GEN_106 = 5'ha == io_ctrl_rs2Addr ? rf__10 : _GEN_105; // @[RegFile.scala 24:{20,20}]
  wire [63:0] _GEN_107 = 5'hb == io_ctrl_rs2Addr ? rf__11 : _GEN_106; // @[RegFile.scala 24:{20,20}]
  wire [63:0] _GEN_108 = 5'hc == io_ctrl_rs2Addr ? rf__12 : _GEN_107; // @[RegFile.scala 24:{20,20}]
  wire [63:0] _GEN_109 = 5'hd == io_ctrl_rs2Addr ? rf__13 : _GEN_108; // @[RegFile.scala 24:{20,20}]
  wire [63:0] _GEN_110 = 5'he == io_ctrl_rs2Addr ? rf__14 : _GEN_109; // @[RegFile.scala 24:{20,20}]
  wire [63:0] _GEN_111 = 5'hf == io_ctrl_rs2Addr ? rf__15 : _GEN_110; // @[RegFile.scala 24:{20,20}]
  wire [63:0] _GEN_112 = 5'h10 == io_ctrl_rs2Addr ? rf__16 : _GEN_111; // @[RegFile.scala 24:{20,20}]
  wire [63:0] _GEN_113 = 5'h11 == io_ctrl_rs2Addr ? rf__17 : _GEN_112; // @[RegFile.scala 24:{20,20}]
  wire [63:0] _GEN_114 = 5'h12 == io_ctrl_rs2Addr ? rf__18 : _GEN_113; // @[RegFile.scala 24:{20,20}]
  wire [63:0] _GEN_115 = 5'h13 == io_ctrl_rs2Addr ? rf__19 : _GEN_114; // @[RegFile.scala 24:{20,20}]
  wire [63:0] _GEN_116 = 5'h14 == io_ctrl_rs2Addr ? rf__20 : _GEN_115; // @[RegFile.scala 24:{20,20}]
  wire [63:0] _GEN_117 = 5'h15 == io_ctrl_rs2Addr ? rf__21 : _GEN_116; // @[RegFile.scala 24:{20,20}]
  wire [63:0] _GEN_118 = 5'h16 == io_ctrl_rs2Addr ? rf__22 : _GEN_117; // @[RegFile.scala 24:{20,20}]
  wire [63:0] _GEN_119 = 5'h17 == io_ctrl_rs2Addr ? rf__23 : _GEN_118; // @[RegFile.scala 24:{20,20}]
  wire [63:0] _GEN_120 = 5'h18 == io_ctrl_rs2Addr ? rf__24 : _GEN_119; // @[RegFile.scala 24:{20,20}]
  wire [63:0] _GEN_121 = 5'h19 == io_ctrl_rs2Addr ? rf__25 : _GEN_120; // @[RegFile.scala 24:{20,20}]
  wire [63:0] _GEN_122 = 5'h1a == io_ctrl_rs2Addr ? rf__26 : _GEN_121; // @[RegFile.scala 24:{20,20}]
  wire [63:0] _GEN_123 = 5'h1b == io_ctrl_rs2Addr ? rf__27 : _GEN_122; // @[RegFile.scala 24:{20,20}]
  wire [63:0] _GEN_124 = 5'h1c == io_ctrl_rs2Addr ? rf__28 : _GEN_123; // @[RegFile.scala 24:{20,20}]
  wire [63:0] _GEN_125 = 5'h1d == io_ctrl_rs2Addr ? rf__29 : _GEN_124; // @[RegFile.scala 24:{20,20}]
  wire [63:0] _GEN_126 = 5'h1e == io_ctrl_rs2Addr ? rf__30 : _GEN_125; // @[RegFile.scala 24:{20,20}]
  wire [63:0] _GEN_127 = 5'h1f == io_ctrl_rs2Addr ? rf__31 : _GEN_126; // @[RegFile.scala 24:{20,20}]
  DifftestArchIntRegState dt_ar ( // @[RegFile.scala 26:21]
    .clock(dt_ar_clock),
    .coreid(dt_ar_coreid),
    .gpr_0(dt_ar_gpr_0),
    .gpr_1(dt_ar_gpr_1),
    .gpr_2(dt_ar_gpr_2),
    .gpr_3(dt_ar_gpr_3),
    .gpr_4(dt_ar_gpr_4),
    .gpr_5(dt_ar_gpr_5),
    .gpr_6(dt_ar_gpr_6),
    .gpr_7(dt_ar_gpr_7),
    .gpr_8(dt_ar_gpr_8),
    .gpr_9(dt_ar_gpr_9),
    .gpr_10(dt_ar_gpr_10),
    .gpr_11(dt_ar_gpr_11),
    .gpr_12(dt_ar_gpr_12),
    .gpr_13(dt_ar_gpr_13),
    .gpr_14(dt_ar_gpr_14),
    .gpr_15(dt_ar_gpr_15),
    .gpr_16(dt_ar_gpr_16),
    .gpr_17(dt_ar_gpr_17),
    .gpr_18(dt_ar_gpr_18),
    .gpr_19(dt_ar_gpr_19),
    .gpr_20(dt_ar_gpr_20),
    .gpr_21(dt_ar_gpr_21),
    .gpr_22(dt_ar_gpr_22),
    .gpr_23(dt_ar_gpr_23),
    .gpr_24(dt_ar_gpr_24),
    .gpr_25(dt_ar_gpr_25),
    .gpr_26(dt_ar_gpr_26),
    .gpr_27(dt_ar_gpr_27),
    .gpr_28(dt_ar_gpr_28),
    .gpr_29(dt_ar_gpr_29),
    .gpr_30(dt_ar_gpr_30),
    .gpr_31(dt_ar_gpr_31)
  );
  assign io_rs1Data = io_ctrl_rs1Addr != 5'h0 & io_ctrl_rs1En ? _GEN_95 : 64'h0; // @[RegFile.scala 23:20]
  assign io_rs2Data = io_ctrl_rs2Addr != 5'h0 & io_ctrl_rs2En ? _GEN_127 : 64'h0; // @[RegFile.scala 24:20]
  assign rf_10 = rf__10;
  assign dt_ar_clock = clock; // @[RegFile.scala 27:19]
  assign dt_ar_coreid = 8'h0; // @[RegFile.scala 28:19]
  assign dt_ar_gpr_0 = rf__0; // @[RegFile.scala 29:19]
  assign dt_ar_gpr_1 = rf__1; // @[RegFile.scala 29:19]
  assign dt_ar_gpr_2 = rf__2; // @[RegFile.scala 29:19]
  assign dt_ar_gpr_3 = rf__3; // @[RegFile.scala 29:19]
  assign dt_ar_gpr_4 = rf__4; // @[RegFile.scala 29:19]
  assign dt_ar_gpr_5 = rf__5; // @[RegFile.scala 29:19]
  assign dt_ar_gpr_6 = rf__6; // @[RegFile.scala 29:19]
  assign dt_ar_gpr_7 = rf__7; // @[RegFile.scala 29:19]
  assign dt_ar_gpr_8 = rf__8; // @[RegFile.scala 29:19]
  assign dt_ar_gpr_9 = rf__9; // @[RegFile.scala 29:19]
  assign dt_ar_gpr_10 = rf__10; // @[RegFile.scala 29:19]
  assign dt_ar_gpr_11 = rf__11; // @[RegFile.scala 29:19]
  assign dt_ar_gpr_12 = rf__12; // @[RegFile.scala 29:19]
  assign dt_ar_gpr_13 = rf__13; // @[RegFile.scala 29:19]
  assign dt_ar_gpr_14 = rf__14; // @[RegFile.scala 29:19]
  assign dt_ar_gpr_15 = rf__15; // @[RegFile.scala 29:19]
  assign dt_ar_gpr_16 = rf__16; // @[RegFile.scala 29:19]
  assign dt_ar_gpr_17 = rf__17; // @[RegFile.scala 29:19]
  assign dt_ar_gpr_18 = rf__18; // @[RegFile.scala 29:19]
  assign dt_ar_gpr_19 = rf__19; // @[RegFile.scala 29:19]
  assign dt_ar_gpr_20 = rf__20; // @[RegFile.scala 29:19]
  assign dt_ar_gpr_21 = rf__21; // @[RegFile.scala 29:19]
  assign dt_ar_gpr_22 = rf__22; // @[RegFile.scala 29:19]
  assign dt_ar_gpr_23 = rf__23; // @[RegFile.scala 29:19]
  assign dt_ar_gpr_24 = rf__24; // @[RegFile.scala 29:19]
  assign dt_ar_gpr_25 = rf__25; // @[RegFile.scala 29:19]
  assign dt_ar_gpr_26 = rf__26; // @[RegFile.scala 29:19]
  assign dt_ar_gpr_27 = rf__27; // @[RegFile.scala 29:19]
  assign dt_ar_gpr_28 = rf__28; // @[RegFile.scala 29:19]
  assign dt_ar_gpr_29 = rf__29; // @[RegFile.scala 29:19]
  assign dt_ar_gpr_30 = rf__30; // @[RegFile.scala 29:19]
  assign dt_ar_gpr_31 = rf__31; // @[RegFile.scala 29:19]
  always @(posedge clock) begin
    if (reset) begin // @[RegFile.scala 17:19]
      rf__0 <= 64'h0; // @[RegFile.scala 17:19]
    end else if (io_rdEn & io_rdAddr != 32'h0) begin // @[RegFile.scala 19:41]
      if (5'h0 == io_rdAddr[4:0]) begin // @[RegFile.scala 20:19]
        rf__0 <= io_rdData; // @[RegFile.scala 20:19]
      end
    end
    if (reset) begin // @[RegFile.scala 17:19]
      rf__1 <= 64'h0; // @[RegFile.scala 17:19]
    end else if (io_rdEn & io_rdAddr != 32'h0) begin // @[RegFile.scala 19:41]
      if (5'h1 == io_rdAddr[4:0]) begin // @[RegFile.scala 20:19]
        rf__1 <= io_rdData; // @[RegFile.scala 20:19]
      end
    end
    if (reset) begin // @[RegFile.scala 17:19]
      rf__2 <= 64'h0; // @[RegFile.scala 17:19]
    end else if (io_rdEn & io_rdAddr != 32'h0) begin // @[RegFile.scala 19:41]
      if (5'h2 == io_rdAddr[4:0]) begin // @[RegFile.scala 20:19]
        rf__2 <= io_rdData; // @[RegFile.scala 20:19]
      end
    end
    if (reset) begin // @[RegFile.scala 17:19]
      rf__3 <= 64'h0; // @[RegFile.scala 17:19]
    end else if (io_rdEn & io_rdAddr != 32'h0) begin // @[RegFile.scala 19:41]
      if (5'h3 == io_rdAddr[4:0]) begin // @[RegFile.scala 20:19]
        rf__3 <= io_rdData; // @[RegFile.scala 20:19]
      end
    end
    if (reset) begin // @[RegFile.scala 17:19]
      rf__4 <= 64'h0; // @[RegFile.scala 17:19]
    end else if (io_rdEn & io_rdAddr != 32'h0) begin // @[RegFile.scala 19:41]
      if (5'h4 == io_rdAddr[4:0]) begin // @[RegFile.scala 20:19]
        rf__4 <= io_rdData; // @[RegFile.scala 20:19]
      end
    end
    if (reset) begin // @[RegFile.scala 17:19]
      rf__5 <= 64'h0; // @[RegFile.scala 17:19]
    end else if (io_rdEn & io_rdAddr != 32'h0) begin // @[RegFile.scala 19:41]
      if (5'h5 == io_rdAddr[4:0]) begin // @[RegFile.scala 20:19]
        rf__5 <= io_rdData; // @[RegFile.scala 20:19]
      end
    end
    if (reset) begin // @[RegFile.scala 17:19]
      rf__6 <= 64'h0; // @[RegFile.scala 17:19]
    end else if (io_rdEn & io_rdAddr != 32'h0) begin // @[RegFile.scala 19:41]
      if (5'h6 == io_rdAddr[4:0]) begin // @[RegFile.scala 20:19]
        rf__6 <= io_rdData; // @[RegFile.scala 20:19]
      end
    end
    if (reset) begin // @[RegFile.scala 17:19]
      rf__7 <= 64'h0; // @[RegFile.scala 17:19]
    end else if (io_rdEn & io_rdAddr != 32'h0) begin // @[RegFile.scala 19:41]
      if (5'h7 == io_rdAddr[4:0]) begin // @[RegFile.scala 20:19]
        rf__7 <= io_rdData; // @[RegFile.scala 20:19]
      end
    end
    if (reset) begin // @[RegFile.scala 17:19]
      rf__8 <= 64'h0; // @[RegFile.scala 17:19]
    end else if (io_rdEn & io_rdAddr != 32'h0) begin // @[RegFile.scala 19:41]
      if (5'h8 == io_rdAddr[4:0]) begin // @[RegFile.scala 20:19]
        rf__8 <= io_rdData; // @[RegFile.scala 20:19]
      end
    end
    if (reset) begin // @[RegFile.scala 17:19]
      rf__9 <= 64'h0; // @[RegFile.scala 17:19]
    end else if (io_rdEn & io_rdAddr != 32'h0) begin // @[RegFile.scala 19:41]
      if (5'h9 == io_rdAddr[4:0]) begin // @[RegFile.scala 20:19]
        rf__9 <= io_rdData; // @[RegFile.scala 20:19]
      end
    end
    if (reset) begin // @[RegFile.scala 17:19]
      rf__10 <= 64'h0; // @[RegFile.scala 17:19]
    end else if (io_rdEn & io_rdAddr != 32'h0) begin // @[RegFile.scala 19:41]
      if (5'ha == io_rdAddr[4:0]) begin // @[RegFile.scala 20:19]
        rf__10 <= io_rdData; // @[RegFile.scala 20:19]
      end
    end
    if (reset) begin // @[RegFile.scala 17:19]
      rf__11 <= 64'h0; // @[RegFile.scala 17:19]
    end else if (io_rdEn & io_rdAddr != 32'h0) begin // @[RegFile.scala 19:41]
      if (5'hb == io_rdAddr[4:0]) begin // @[RegFile.scala 20:19]
        rf__11 <= io_rdData; // @[RegFile.scala 20:19]
      end
    end
    if (reset) begin // @[RegFile.scala 17:19]
      rf__12 <= 64'h0; // @[RegFile.scala 17:19]
    end else if (io_rdEn & io_rdAddr != 32'h0) begin // @[RegFile.scala 19:41]
      if (5'hc == io_rdAddr[4:0]) begin // @[RegFile.scala 20:19]
        rf__12 <= io_rdData; // @[RegFile.scala 20:19]
      end
    end
    if (reset) begin // @[RegFile.scala 17:19]
      rf__13 <= 64'h0; // @[RegFile.scala 17:19]
    end else if (io_rdEn & io_rdAddr != 32'h0) begin // @[RegFile.scala 19:41]
      if (5'hd == io_rdAddr[4:0]) begin // @[RegFile.scala 20:19]
        rf__13 <= io_rdData; // @[RegFile.scala 20:19]
      end
    end
    if (reset) begin // @[RegFile.scala 17:19]
      rf__14 <= 64'h0; // @[RegFile.scala 17:19]
    end else if (io_rdEn & io_rdAddr != 32'h0) begin // @[RegFile.scala 19:41]
      if (5'he == io_rdAddr[4:0]) begin // @[RegFile.scala 20:19]
        rf__14 <= io_rdData; // @[RegFile.scala 20:19]
      end
    end
    if (reset) begin // @[RegFile.scala 17:19]
      rf__15 <= 64'h0; // @[RegFile.scala 17:19]
    end else if (io_rdEn & io_rdAddr != 32'h0) begin // @[RegFile.scala 19:41]
      if (5'hf == io_rdAddr[4:0]) begin // @[RegFile.scala 20:19]
        rf__15 <= io_rdData; // @[RegFile.scala 20:19]
      end
    end
    if (reset) begin // @[RegFile.scala 17:19]
      rf__16 <= 64'h0; // @[RegFile.scala 17:19]
    end else if (io_rdEn & io_rdAddr != 32'h0) begin // @[RegFile.scala 19:41]
      if (5'h10 == io_rdAddr[4:0]) begin // @[RegFile.scala 20:19]
        rf__16 <= io_rdData; // @[RegFile.scala 20:19]
      end
    end
    if (reset) begin // @[RegFile.scala 17:19]
      rf__17 <= 64'h0; // @[RegFile.scala 17:19]
    end else if (io_rdEn & io_rdAddr != 32'h0) begin // @[RegFile.scala 19:41]
      if (5'h11 == io_rdAddr[4:0]) begin // @[RegFile.scala 20:19]
        rf__17 <= io_rdData; // @[RegFile.scala 20:19]
      end
    end
    if (reset) begin // @[RegFile.scala 17:19]
      rf__18 <= 64'h0; // @[RegFile.scala 17:19]
    end else if (io_rdEn & io_rdAddr != 32'h0) begin // @[RegFile.scala 19:41]
      if (5'h12 == io_rdAddr[4:0]) begin // @[RegFile.scala 20:19]
        rf__18 <= io_rdData; // @[RegFile.scala 20:19]
      end
    end
    if (reset) begin // @[RegFile.scala 17:19]
      rf__19 <= 64'h0; // @[RegFile.scala 17:19]
    end else if (io_rdEn & io_rdAddr != 32'h0) begin // @[RegFile.scala 19:41]
      if (5'h13 == io_rdAddr[4:0]) begin // @[RegFile.scala 20:19]
        rf__19 <= io_rdData; // @[RegFile.scala 20:19]
      end
    end
    if (reset) begin // @[RegFile.scala 17:19]
      rf__20 <= 64'h0; // @[RegFile.scala 17:19]
    end else if (io_rdEn & io_rdAddr != 32'h0) begin // @[RegFile.scala 19:41]
      if (5'h14 == io_rdAddr[4:0]) begin // @[RegFile.scala 20:19]
        rf__20 <= io_rdData; // @[RegFile.scala 20:19]
      end
    end
    if (reset) begin // @[RegFile.scala 17:19]
      rf__21 <= 64'h0; // @[RegFile.scala 17:19]
    end else if (io_rdEn & io_rdAddr != 32'h0) begin // @[RegFile.scala 19:41]
      if (5'h15 == io_rdAddr[4:0]) begin // @[RegFile.scala 20:19]
        rf__21 <= io_rdData; // @[RegFile.scala 20:19]
      end
    end
    if (reset) begin // @[RegFile.scala 17:19]
      rf__22 <= 64'h0; // @[RegFile.scala 17:19]
    end else if (io_rdEn & io_rdAddr != 32'h0) begin // @[RegFile.scala 19:41]
      if (5'h16 == io_rdAddr[4:0]) begin // @[RegFile.scala 20:19]
        rf__22 <= io_rdData; // @[RegFile.scala 20:19]
      end
    end
    if (reset) begin // @[RegFile.scala 17:19]
      rf__23 <= 64'h0; // @[RegFile.scala 17:19]
    end else if (io_rdEn & io_rdAddr != 32'h0) begin // @[RegFile.scala 19:41]
      if (5'h17 == io_rdAddr[4:0]) begin // @[RegFile.scala 20:19]
        rf__23 <= io_rdData; // @[RegFile.scala 20:19]
      end
    end
    if (reset) begin // @[RegFile.scala 17:19]
      rf__24 <= 64'h0; // @[RegFile.scala 17:19]
    end else if (io_rdEn & io_rdAddr != 32'h0) begin // @[RegFile.scala 19:41]
      if (5'h18 == io_rdAddr[4:0]) begin // @[RegFile.scala 20:19]
        rf__24 <= io_rdData; // @[RegFile.scala 20:19]
      end
    end
    if (reset) begin // @[RegFile.scala 17:19]
      rf__25 <= 64'h0; // @[RegFile.scala 17:19]
    end else if (io_rdEn & io_rdAddr != 32'h0) begin // @[RegFile.scala 19:41]
      if (5'h19 == io_rdAddr[4:0]) begin // @[RegFile.scala 20:19]
        rf__25 <= io_rdData; // @[RegFile.scala 20:19]
      end
    end
    if (reset) begin // @[RegFile.scala 17:19]
      rf__26 <= 64'h0; // @[RegFile.scala 17:19]
    end else if (io_rdEn & io_rdAddr != 32'h0) begin // @[RegFile.scala 19:41]
      if (5'h1a == io_rdAddr[4:0]) begin // @[RegFile.scala 20:19]
        rf__26 <= io_rdData; // @[RegFile.scala 20:19]
      end
    end
    if (reset) begin // @[RegFile.scala 17:19]
      rf__27 <= 64'h0; // @[RegFile.scala 17:19]
    end else if (io_rdEn & io_rdAddr != 32'h0) begin // @[RegFile.scala 19:41]
      if (5'h1b == io_rdAddr[4:0]) begin // @[RegFile.scala 20:19]
        rf__27 <= io_rdData; // @[RegFile.scala 20:19]
      end
    end
    if (reset) begin // @[RegFile.scala 17:19]
      rf__28 <= 64'h0; // @[RegFile.scala 17:19]
    end else if (io_rdEn & io_rdAddr != 32'h0) begin // @[RegFile.scala 19:41]
      if (5'h1c == io_rdAddr[4:0]) begin // @[RegFile.scala 20:19]
        rf__28 <= io_rdData; // @[RegFile.scala 20:19]
      end
    end
    if (reset) begin // @[RegFile.scala 17:19]
      rf__29 <= 64'h0; // @[RegFile.scala 17:19]
    end else if (io_rdEn & io_rdAddr != 32'h0) begin // @[RegFile.scala 19:41]
      if (5'h1d == io_rdAddr[4:0]) begin // @[RegFile.scala 20:19]
        rf__29 <= io_rdData; // @[RegFile.scala 20:19]
      end
    end
    if (reset) begin // @[RegFile.scala 17:19]
      rf__30 <= 64'h0; // @[RegFile.scala 17:19]
    end else if (io_rdEn & io_rdAddr != 32'h0) begin // @[RegFile.scala 19:41]
      if (5'h1e == io_rdAddr[4:0]) begin // @[RegFile.scala 20:19]
        rf__30 <= io_rdData; // @[RegFile.scala 20:19]
      end
    end
    if (reset) begin // @[RegFile.scala 17:19]
      rf__31 <= 64'h0; // @[RegFile.scala 17:19]
    end else if (io_rdEn & io_rdAddr != 32'h0) begin // @[RegFile.scala 19:41]
      if (5'h1f == io_rdAddr[4:0]) begin // @[RegFile.scala 20:19]
        rf__31 <= io_rdData; // @[RegFile.scala 20:19]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  rf__0 = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  rf__1 = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  rf__2 = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  rf__3 = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  rf__4 = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  rf__5 = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  rf__6 = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  rf__7 = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  rf__8 = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  rf__9 = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  rf__10 = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  rf__11 = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  rf__12 = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  rf__13 = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  rf__14 = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  rf__15 = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  rf__16 = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  rf__17 = _RAND_17[63:0];
  _RAND_18 = {2{`RANDOM}};
  rf__18 = _RAND_18[63:0];
  _RAND_19 = {2{`RANDOM}};
  rf__19 = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  rf__20 = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  rf__21 = _RAND_21[63:0];
  _RAND_22 = {2{`RANDOM}};
  rf__22 = _RAND_22[63:0];
  _RAND_23 = {2{`RANDOM}};
  rf__23 = _RAND_23[63:0];
  _RAND_24 = {2{`RANDOM}};
  rf__24 = _RAND_24[63:0];
  _RAND_25 = {2{`RANDOM}};
  rf__25 = _RAND_25[63:0];
  _RAND_26 = {2{`RANDOM}};
  rf__26 = _RAND_26[63:0];
  _RAND_27 = {2{`RANDOM}};
  rf__27 = _RAND_27[63:0];
  _RAND_28 = {2{`RANDOM}};
  rf__28 = _RAND_28[63:0];
  _RAND_29 = {2{`RANDOM}};
  rf__29 = _RAND_29[63:0];
  _RAND_30 = {2{`RANDOM}};
  rf__30 = _RAND_30[63:0];
  _RAND_31 = {2{`RANDOM}};
  rf__31 = _RAND_31[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ImmGen(
  input  [31:0] io_inst,
  input  [2:0]  io_immOp,
  output [63:0] io_imm
);
  wire [51:0] _immType_0_T_2 = io_inst[31] ? 52'hfffffffffffff : 52'h0; // @[Bitwise.scala 74:12]
  wire [63:0] immType_0 = {_immType_0_T_2,io_inst[31:20]}; // @[ImmGen.scala 19:41]
  wire [31:0] _immType_1_T_2 = io_inst[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] immType_1 = {_immType_1_T_2,io_inst[31:12],12'h0}; // @[ImmGen.scala 20:59]
  wire [63:0] immType_2 = {_immType_0_T_2,io_inst[31:25],io_inst[11:7]}; // @[ImmGen.scala 21:59]
  wire [64:0] _immType_3_T_11 = {_immType_0_T_2,io_inst[31],io_inst[7],io_inst[30:25],io_inst[11:8],1'h0}; // @[ImmGen.scala 22:113]
  wire [42:0] _immType_4_T_2 = io_inst[31] ? 43'h7ffffffffff : 43'h0; // @[Bitwise.scala 74:12]
  wire [63:0] immType_4 = {_immType_4_T_2,io_inst[31],io_inst[19:12],io_inst[20],io_inst[30:21],1'h0}; // @[ImmGen.scala 23:113]
  wire [63:0] _GEN_1 = 3'h1 == io_immOp ? immType_1 : immType_0; // @[ImmGen.scala 25:{10,10}]
  wire [63:0] _GEN_2 = 3'h2 == io_immOp ? immType_2 : _GEN_1; // @[ImmGen.scala 25:{10,10}]
  wire [63:0] immType_3 = _immType_3_T_11[63:0]; // @[ImmGen.scala 17:21 22:16]
  wire [63:0] _GEN_3 = 3'h3 == io_immOp ? immType_3 : _GEN_2; // @[ImmGen.scala 25:{10,10}]
  assign io_imm = 3'h4 == io_immOp ? immType_4 : _GEN_3; // @[ImmGen.scala 25:{10,10}]
endmodule
module ContrGen(
  input  [31:0] io_inst,
  output [2:0]  io_branch,
  output [2:0]  io_immOp,
  output        io_rdEn,
  output [4:0]  io_rdAddr,
  output        io_typeL,
  output        io_aluCtr_aluA,
  output [1:0]  io_aluCtr_aluB,
  output [3:0]  io_aluCtr_aluOp,
  output [1:0]  io_memCtr_memtoReg,
  output        io_memCtr_memWr,
  output [2:0]  io_memCtr_memOP,
  output        io_regCtrl_rs1En,
  output        io_regCtrl_rs2En,
  output [4:0]  io_regCtrl_rs1Addr,
  output [4:0]  io_regCtrl_rs2Addr
);
  wire [31:0] _instLui_T = io_inst & 32'h7f; // @[ContrGen.scala 24:26]
  wire  instLui = 32'h37 == _instLui_T; // @[ContrGen.scala 24:26]
  wire  instAuipc = 32'h17 == _instLui_T; // @[ContrGen.scala 25:26]
  wire  typeU = instLui | instAuipc; // @[ContrGen.scala 26:29]
  wire [31:0] _instAddi_T = io_inst & 32'h707f; // @[ContrGen.scala 28:26]
  wire  instAddi = 32'h13 == _instAddi_T; // @[ContrGen.scala 28:26]
  wire  instAndi = 32'h7013 == _instAddi_T; // @[ContrGen.scala 29:26]
  wire  instXori = 32'h4013 == _instAddi_T; // @[ContrGen.scala 30:26]
  wire  instOri = 32'h6013 == _instAddi_T; // @[ContrGen.scala 31:26]
  wire [31:0] _instSlli_T = io_inst & 32'hfc00707f; // @[ContrGen.scala 32:26]
  wire  instSlli = 32'h1013 == _instSlli_T; // @[ContrGen.scala 32:26]
  wire  instSrli = 32'h5013 == _instSlli_T; // @[ContrGen.scala 33:26]
  wire  instSrai = 32'h40005013 == _instSlli_T; // @[ContrGen.scala 34:26]
  wire  instSlti = 32'h2013 == _instAddi_T; // @[ContrGen.scala 35:26]
  wire  instSltiu = 32'h3013 == _instAddi_T; // @[ContrGen.scala 36:26]
  wire  instAddiw = 32'h1b == _instAddi_T; // @[ContrGen.scala 37:26]
  wire [31:0] _instSlliw_T = io_inst & 32'hfe00707f; // @[ContrGen.scala 38:26]
  wire  instSlliw = 32'h101b == _instSlliw_T; // @[ContrGen.scala 38:26]
  wire  instSrliw = 32'h501b == _instSlliw_T; // @[ContrGen.scala 39:26]
  wire  instSraiw = 32'h4000501b == _instSlliw_T; // @[ContrGen.scala 40:26]
  wire  instJalr = 32'h67 == _instAddi_T; // @[ContrGen.scala 41:26]
  wire  instLb = 32'h3 == _instAddi_T; // @[ContrGen.scala 42:26]
  wire  instLh = 32'h1003 == _instAddi_T; // @[ContrGen.scala 43:26]
  wire  instLw = 32'h2003 == _instAddi_T; // @[ContrGen.scala 44:26]
  wire  instLd = 32'h3003 == _instAddi_T; // @[ContrGen.scala 45:26]
  wire  instLbu = 32'h4003 == _instAddi_T; // @[ContrGen.scala 46:26]
  wire  instLhu = 32'h5003 == _instAddi_T; // @[ContrGen.scala 47:26]
  wire  instLwu = 32'h6003 == _instAddi_T; // @[ContrGen.scala 48:26]
  wire  _typeL_T_1 = instLb | instLh | instLw; // @[ContrGen.scala 53:32]
  wire  _typeL_T_4 = instLb | instLh | instLw | instLd | instLbu | instLhu; // @[ContrGen.scala 53:63]
  wire  instJal = 32'h6f == _instLui_T; // @[ContrGen.scala 56:26]
  wire  typeJ = instJal | instJalr; // @[ContrGen.scala 57:29]
  wire  instAdd = 32'h33 == _instSlliw_T; // @[ContrGen.scala 59:26]
  wire  instSub = 32'h40000033 == _instSlliw_T; // @[ContrGen.scala 60:26]
  wire  instSll = 32'h1033 == _instSlliw_T; // @[ContrGen.scala 61:26]
  wire  instSlt = 32'h2033 == _instSlliw_T; // @[ContrGen.scala 62:26]
  wire  instSltu = 32'h3033 == _instSlliw_T; // @[ContrGen.scala 63:26]
  wire  instXor = 32'h4033 == _instSlliw_T; // @[ContrGen.scala 64:26]
  wire  instSrl = 32'h5033 == _instSlliw_T; // @[ContrGen.scala 65:26]
  wire  instSra = 32'h40005033 == _instSlliw_T; // @[ContrGen.scala 66:26]
  wire  instOr = 32'h6033 == _instSlliw_T; // @[ContrGen.scala 67:26]
  wire  instAnd = 32'h7033 == _instSlliw_T; // @[ContrGen.scala 68:26]
  wire  instAddw = 32'h3b == _instSlliw_T; // @[ContrGen.scala 69:26]
  wire  instSubw = 32'h4000003b == _instSlliw_T; // @[ContrGen.scala 70:26]
  wire  instSllw = 32'h103b == _instSlliw_T; // @[ContrGen.scala 71:26]
  wire  instSrlw = 32'h503b == _instSlliw_T; // @[ContrGen.scala 72:26]
  wire  instSraw = 32'h4000503b == _instSlliw_T; // @[ContrGen.scala 73:26]
  wire  instMret = 32'h30200073 == io_inst; // @[ContrGen.scala 74:26]
  wire  aluRem = 32'h200603b == _instSlliw_T; // @[ContrGen.scala 75:26]
  wire  instDiv = 32'h2004033 == _instSlliw_T; // @[ContrGen.scala 76:26]
  wire  instDivw = 32'h200403b == _instSlliw_T; // @[ContrGen.scala 77:26]
  wire  instMul = 32'h2000033 == _instSlliw_T; // @[ContrGen.scala 78:26]
  wire  instMulw = 32'h200003b == _instSlliw_T; // @[ContrGen.scala 79:26]
  wire  _typeR_T_4 = instAdd | instSub | instSll | instSlt | instSltu | instXor; // @[ContrGen.scala 80:78]
  wire  _typeR_T_9 = _typeR_T_4 | instSrl | instSra | instOr | instAnd | instAddw; // @[ContrGen.scala 81:78]
  wire  _typeR_T_14 = _typeR_T_9 | instSubw | instSllw | instSrlw | instSraw | instMret; // @[ContrGen.scala 82:78]
  wire  typeR = _typeR_T_14 | aluRem | instDiv | instDivw | instMul | instMulw; // @[ContrGen.scala 83:78]
  wire  instBeq = 32'h63 == _instAddi_T; // @[ContrGen.scala 85:27]
  wire  instBne = 32'h1063 == _instAddi_T; // @[ContrGen.scala 86:27]
  wire  instBlt = 32'h4063 == _instAddi_T; // @[ContrGen.scala 87:27]
  wire  instBge = 32'h5063 == _instAddi_T; // @[ContrGen.scala 88:27]
  wire  instBltu = 32'h6063 == _instAddi_T; // @[ContrGen.scala 89:27]
  wire  instBgeu = 32'h7063 == _instAddi_T; // @[ContrGen.scala 90:27]
  wire  _typeB_T = instBeq | instBne; // @[ContrGen.scala 91:30]
  wire  typeB = instBeq | instBne | instBlt | instBge | instBltu | instBgeu; // @[ContrGen.scala 91:74]
  wire  instSb = 32'h23 == _instAddi_T; // @[ContrGen.scala 93:27]
  wire  instSh = 32'h1023 == _instAddi_T; // @[ContrGen.scala 94:27]
  wire  instSw = 32'h2023 == _instAddi_T; // @[ContrGen.scala 95:27]
  wire  instSd = 32'h3023 == _instAddi_T; // @[ContrGen.scala 96:27]
  wire  _typeS_T_1 = instSb | instSh | instSw; // @[ContrGen.scala 97:39]
  wire  typeS = instSb | instSh | instSw | instSd; // @[ContrGen.scala 97:49]
  wire  Ebreak = 32'h100073 == io_inst; // @[ContrGen.scala 99:27]
  wire  _typeW_T_3 = instAddw | instSubw | instSllw | instSlliw | instSraw; // @[ContrGen.scala 101:68]
  wire  _typeW_T_9 = _typeW_T_3 | instSrlw | instSrliw | instSraiw | instAddiw | aluRem | instDivw; // @[ContrGen.scala 102:76]
  wire  typeW = _typeW_T_9 | instMulw; // @[ContrGen.scala 103:14]
  wire  _io_aluCtr_aluB_T = typeR | typeB; // @[ContrGen.scala 109:12]
  wire [1:0] _io_aluCtr_aluB_T_1 = typeJ ? 2'h2 : 2'h1; // @[Mux.scala 101:16]
  wire  aluSub = instSub | instSubw; // @[ContrGen.scala 116:28]
  wire  aluSlt = instSlti | instSlt; // @[ContrGen.scala 117:29]
  wire  aluSltu = instSltiu | instSltu; // @[ContrGen.scala 118:29]
  wire  aluAnd = instAndi | instAnd; // @[ContrGen.scala 119:29]
  wire  aluOr = instOri | instOr; // @[ContrGen.scala 120:29]
  wire  aluXor = instXori | instXor; // @[ContrGen.scala 121:29]
  wire  aluSll = instSlli | instSlliw | instSll | instSllw; // @[ContrGen.scala 122:53]
  wire  aluSrl = instSrli | instSrliw | instSrl | instSrlw; // @[ContrGen.scala 123:53]
  wire  aluSra = instSrai | instSraiw | instSra | instSraw; // @[ContrGen.scala 124:53]
  wire  aluDiv = instDiv | instDivw; // @[ContrGen.scala 126:27]
  wire  aluMul = instMul | instMulw; // @[ContrGen.scala 127:27]
  wire  _io_aluCtr_aluOp_T_2 = aluSlt | instBlt | instBge; // @[ContrGen.scala 133:37]
  wire  _io_aluCtr_aluOp_T_6 = aluSltu | instBltu | instBgeu; // @[ContrGen.scala 135:40]
  wire [2:0] _io_aluCtr_aluOp_T_7 = aluAnd ? 3'h7 : 3'h0; // @[Mux.scala 101:16]
  wire [3:0] _io_aluCtr_aluOp_T_8 = aluMul ? 4'he : {{1'd0}, _io_aluCtr_aluOp_T_7}; // @[Mux.scala 101:16]
  wire [3:0] _io_aluCtr_aluOp_T_9 = aluOr ? 4'h6 : _io_aluCtr_aluOp_T_8; // @[Mux.scala 101:16]
  wire [3:0] _io_aluCtr_aluOp_T_10 = aluSra ? 4'hd : _io_aluCtr_aluOp_T_9; // @[Mux.scala 101:16]
  wire [3:0] _io_aluCtr_aluOp_T_11 = aluSrl ? 4'h5 : _io_aluCtr_aluOp_T_10; // @[Mux.scala 101:16]
  wire [3:0] _io_aluCtr_aluOp_T_12 = aluDiv ? 4'hc : _io_aluCtr_aluOp_T_11; // @[Mux.scala 101:16]
  wire [3:0] _io_aluCtr_aluOp_T_13 = aluXor ? 4'h4 : _io_aluCtr_aluOp_T_12; // @[Mux.scala 101:16]
  wire [3:0] _io_aluCtr_aluOp_T_14 = aluRem ? 4'hb : _io_aluCtr_aluOp_T_13; // @[Mux.scala 101:16]
  wire [3:0] _io_aluCtr_aluOp_T_15 = instLui ? 4'h3 : _io_aluCtr_aluOp_T_14; // @[Mux.scala 101:16]
  wire [3:0] _io_aluCtr_aluOp_T_16 = _io_aluCtr_aluOp_T_6 ? 4'ha : _io_aluCtr_aluOp_T_15; // @[Mux.scala 101:16]
  wire [3:0] _io_aluCtr_aluOp_T_17 = _typeB_T ? 4'h9 : _io_aluCtr_aluOp_T_16; // @[Mux.scala 101:16]
  wire [3:0] _io_aluCtr_aluOp_T_18 = _io_aluCtr_aluOp_T_2 ? 4'h2 : _io_aluCtr_aluOp_T_17; // @[Mux.scala 101:16]
  wire [3:0] _io_aluCtr_aluOp_T_19 = aluSll ? 4'h1 : _io_aluCtr_aluOp_T_18; // @[Mux.scala 101:16]
  wire  _io_branch_T = instBlt | instBltu; // @[ContrGen.scala 151:20]
  wire  _io_branch_T_1 = instBge | instBgeu; // @[ContrGen.scala 152:20]
  wire [2:0] _io_branch_T_2 = _io_branch_T_1 ? 3'h7 : 3'h0; // @[Mux.scala 101:16]
  wire [2:0] _io_branch_T_3 = _io_branch_T ? 3'h6 : _io_branch_T_2; // @[Mux.scala 101:16]
  wire [2:0] _io_branch_T_4 = instBne ? 3'h5 : _io_branch_T_3; // @[Mux.scala 101:16]
  wire [2:0] _io_branch_T_5 = instBeq ? 3'h4 : _io_branch_T_4; // @[Mux.scala 101:16]
  wire [2:0] _io_branch_T_6 = instJalr ? 3'h2 : _io_branch_T_5; // @[Mux.scala 101:16]
  wire  wRegEn = ~(typeS | typeB | Ebreak); // @[ContrGen.scala 159:16]
  wire  _io_immOp_T_8 = instAddi | instAddiw | instSlti | instSltiu | instXori | instOri | instAndi | instSlli |
    instSlliw | instSrli; // @[ContrGen.scala 164:120]
  wire  _io_immOp_T_15 = _io_immOp_T_8 | instSrliw | instSrai | instSraiw | instJalr | instLb | instLh | instLw; // @[ContrGen.scala 165:92]
  wire  _io_immOp_T_19 = _io_immOp_T_15 | instLwu | instLd | instLbu | instLhu; // @[ContrGen.scala 166:57]
  wire  _io_immOp_T_20 = instAuipc | instLui; // @[ContrGen.scala 167:22]
  wire  _io_immOp_T_23 = instSd | instSb | instSw | instSh; // @[ContrGen.scala 168:39]
  wire [2:0] _io_immOp_T_29 = instJal ? 3'h4 : 3'h7; // @[Mux.scala 101:16]
  wire [2:0] _io_immOp_T_30 = typeB ? 3'h3 : _io_immOp_T_29; // @[Mux.scala 101:16]
  wire [2:0] _io_immOp_T_31 = _io_immOp_T_23 ? 3'h2 : _io_immOp_T_30; // @[Mux.scala 101:16]
  wire [2:0] _io_immOp_T_32 = _io_immOp_T_20 ? 3'h1 : _io_immOp_T_31; // @[Mux.scala 101:16]
  wire  _io_memCtr_memtoReg_T_5 = _typeL_T_1 | instLwu | instLd | instLbu | instLhu; // @[ContrGen.scala 173:65]
  wire [1:0] _io_memCtr_memtoReg_T_6 = typeW ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire  _io_memCtr_memOP_T = instLb | instSb; // @[ContrGen.scala 179:19]
  wire  _io_memCtr_memOP_T_1 = instLh | instSh; // @[ContrGen.scala 180:19]
  wire  _io_memCtr_memOP_T_2 = instLw | instSw; // @[ContrGen.scala 181:19]
  wire  _io_memCtr_memOP_T_3 = instLd | instSd; // @[ContrGen.scala 182:19]
  wire [2:0] _io_memCtr_memOP_T_4 = instLwu ? 3'h6 : 3'h7; // @[Mux.scala 101:16]
  wire [2:0] _io_memCtr_memOP_T_5 = instLhu ? 3'h5 : _io_memCtr_memOP_T_4; // @[Mux.scala 101:16]
  wire [2:0] _io_memCtr_memOP_T_6 = instLbu ? 3'h4 : _io_memCtr_memOP_T_5; // @[Mux.scala 101:16]
  wire [2:0] _io_memCtr_memOP_T_7 = _io_memCtr_memOP_T_3 ? 3'h3 : _io_memCtr_memOP_T_6; // @[Mux.scala 101:16]
  wire [2:0] _io_memCtr_memOP_T_8 = _io_memCtr_memOP_T_2 ? 3'h2 : _io_memCtr_memOP_T_7; // @[Mux.scala 101:16]
  wire [2:0] _io_memCtr_memOP_T_9 = _io_memCtr_memOP_T_1 ? 3'h1 : _io_memCtr_memOP_T_8; // @[Mux.scala 101:16]
  assign io_branch = instJal ? 3'h1 : _io_branch_T_6; // @[Mux.scala 101:16]
  assign io_immOp = _io_immOp_T_19 ? 3'h0 : _io_immOp_T_32; // @[Mux.scala 101:16]
  assign io_rdEn = ~(typeS | typeB | Ebreak); // @[ContrGen.scala 159:16]
  assign io_rdAddr = wRegEn ? io_inst[11:7] : 5'h0; // @[ContrGen.scala 161:19]
  assign io_typeL = _typeL_T_4 | instLwu; // @[ContrGen.scala 54:22]
  assign io_aluCtr_aluA = instAuipc | typeJ; // @[ContrGen.scala 106:35]
  assign io_aluCtr_aluB = _io_aluCtr_aluB_T ? 2'h0 : _io_aluCtr_aluB_T_1; // @[Mux.scala 101:16]
  assign io_aluCtr_aluOp = aluSub ? 4'h8 : _io_aluCtr_aluOp_T_19; // @[Mux.scala 101:16]
  assign io_memCtr_memtoReg = _io_memCtr_memtoReg_T_5 ? 2'h1 : _io_memCtr_memtoReg_T_6; // @[Mux.scala 101:16]
  assign io_memCtr_memWr = _typeS_T_1 | instSd; // @[ContrGen.scala 177:56]
  assign io_memCtr_memOP = _io_memCtr_memOP_T ? 3'h0 : _io_memCtr_memOP_T_9; // @[Mux.scala 101:16]
  assign io_regCtrl_rs1En = ~(typeU | instJal); // @[ContrGen.scala 154:23]
  assign io_regCtrl_rs2En = _io_aluCtr_aluB_T | typeS; // @[ContrGen.scala 155:40]
  assign io_regCtrl_rs1Addr = Ebreak ? 5'ha : io_inst[19:15]; // @[ContrGen.scala 156:28]
  assign io_regCtrl_rs2Addr = io_inst[24:20]; // @[ContrGen.scala 157:29]
endmodule
module Decode(
  input         clock,
  input         reset,
  input         io_rdEn,
  input  [4:0]  io_rdAddr,
  input  [63:0] io_rdData,
  input         io_in_valid,
  input  [31:0] io_in_pc,
  input  [31:0] io_in_inst,
  input         io_exeRdEn,
  input  [4:0]  io_exeRdAddr,
  input  [63:0] io_exeRdData,
  input         io_memRdEn,
  input  [4:0]  io_memRdAddr,
  input  [63:0] io_memRdData,
  input         io_wbRdEn,
  input  [4:0]  io_wbRdAddr,
  input  [63:0] io_wbRdData,
  output        io_bubbleId,
  output        io_out_valid,
  output [31:0] io_out_pc,
  output [31:0] io_out_inst,
  output        io_out_typeL,
  output        io_out_aluA,
  output [1:0]  io_out_aluB,
  output [3:0]  io_out_aluOp,
  output [2:0]  io_out_branch,
  output [1:0]  io_out_memtoReg,
  output        io_out_memWr,
  output [2:0]  io_out_memOp,
  output        io_out_rdEn,
  output [4:0]  io_out_rdAddr,
  output [63:0] io_out_rs1Data,
  output [63:0] io_out_rs2Data,
  output [63:0] io_out_imm,
  output [63:0] rf_10
);
  wire  regs_clock; // @[Decode.scala 35:20]
  wire  regs_reset; // @[Decode.scala 35:20]
  wire [63:0] regs_io_rs1Data; // @[Decode.scala 35:20]
  wire [63:0] regs_io_rs2Data; // @[Decode.scala 35:20]
  wire  regs_io_rdEn; // @[Decode.scala 35:20]
  wire [31:0] regs_io_rdAddr; // @[Decode.scala 35:20]
  wire [63:0] regs_io_rdData; // @[Decode.scala 35:20]
  wire  regs_io_ctrl_rs1En; // @[Decode.scala 35:20]
  wire  regs_io_ctrl_rs2En; // @[Decode.scala 35:20]
  wire [4:0] regs_io_ctrl_rs1Addr; // @[Decode.scala 35:20]
  wire [4:0] regs_io_ctrl_rs2Addr; // @[Decode.scala 35:20]
  wire [63:0] regs_rf_10; // @[Decode.scala 35:20]
  wire [31:0] imm_io_inst; // @[Decode.scala 36:20]
  wire [2:0] imm_io_immOp; // @[Decode.scala 36:20]
  wire [63:0] imm_io_imm; // @[Decode.scala 36:20]
  wire [31:0] con_io_inst; // @[Decode.scala 37:20]
  wire [2:0] con_io_branch; // @[Decode.scala 37:20]
  wire [2:0] con_io_immOp; // @[Decode.scala 37:20]
  wire  con_io_rdEn; // @[Decode.scala 37:20]
  wire [4:0] con_io_rdAddr; // @[Decode.scala 37:20]
  wire  con_io_typeL; // @[Decode.scala 37:20]
  wire  con_io_aluCtr_aluA; // @[Decode.scala 37:20]
  wire [1:0] con_io_aluCtr_aluB; // @[Decode.scala 37:20]
  wire [3:0] con_io_aluCtr_aluOp; // @[Decode.scala 37:20]
  wire [1:0] con_io_memCtr_memtoReg; // @[Decode.scala 37:20]
  wire  con_io_memCtr_memWr; // @[Decode.scala 37:20]
  wire [2:0] con_io_memCtr_memOP; // @[Decode.scala 37:20]
  wire  con_io_regCtrl_rs1En; // @[Decode.scala 37:20]
  wire  con_io_regCtrl_rs2En; // @[Decode.scala 37:20]
  wire [4:0] con_io_regCtrl_rs1Addr; // @[Decode.scala 37:20]
  wire [4:0] con_io_regCtrl_rs2Addr; // @[Decode.scala 37:20]
  wire [4:0] rs1Addr = con_io_regCtrl_rs1En ? con_io_regCtrl_rs1Addr : 5'h0; // @[Decode.scala 50:20]
  wire [4:0] rs2Addr = con_io_regCtrl_rs2En ? con_io_regCtrl_rs2Addr : 5'h0; // @[Decode.scala 51:20]
  wire  _rdRs1HitEx_T_2 = rs1Addr != 5'h0; // @[Decode.scala 52:73]
  wire  rdRs1HitEx = io_exeRdEn & rs1Addr == io_exeRdAddr & rs1Addr != 5'h0; // @[Decode.scala 52:61]
  wire  rdRs1HitMem = io_memRdEn & rs1Addr == io_memRdAddr & _rdRs1HitEx_T_2; // @[Decode.scala 53:62]
  wire  rdRs1HitWb = io_wbRdEn & rs1Addr == io_wbRdAddr & _rdRs1HitEx_T_2; // @[Decode.scala 54:59]
  wire  _rdRs2HitEx_T_2 = rs2Addr != 5'h0; // @[Decode.scala 56:73]
  wire  rdRs2HitEx = io_exeRdEn & rs2Addr == io_exeRdAddr & rs2Addr != 5'h0; // @[Decode.scala 56:61]
  wire  rdRs2HitMem = io_memRdEn & rs2Addr == io_memRdAddr & _rdRs2HitEx_T_2; // @[Decode.scala 57:62]
  wire  rdRs2HitWb = io_wbRdEn & rs2Addr == io_wbRdAddr & _rdRs2HitEx_T_2; // @[Decode.scala 58:59]
  wire [63:0] _rs1Data_T = rdRs1HitWb ? io_wbRdData : regs_io_rs1Data; // @[Decode.scala 63:8]
  wire [63:0] _rs1Data_T_1 = rdRs1HitMem ? io_memRdData : _rs1Data_T; // @[Decode.scala 62:8]
  wire [63:0] _rs1Data_T_2 = rdRs1HitEx ? io_exeRdData : _rs1Data_T_1; // @[Decode.scala 61:8]
  wire [63:0] _rs2Data_T = rdRs2HitWb ? io_wbRdData : regs_io_rs2Data; // @[Decode.scala 68:8]
  wire [63:0] _rs2Data_T_1 = rdRs2HitMem ? io_memRdData : _rs2Data_T; // @[Decode.scala 67:8]
  wire [63:0] _rs2Data_T_2 = rdRs2HitEx ? io_exeRdData : _rs2Data_T_1; // @[Decode.scala 66:8]
  RegFile regs ( // @[Decode.scala 35:20]
    .clock(regs_clock),
    .reset(regs_reset),
    .io_rs1Data(regs_io_rs1Data),
    .io_rs2Data(regs_io_rs2Data),
    .io_rdEn(regs_io_rdEn),
    .io_rdAddr(regs_io_rdAddr),
    .io_rdData(regs_io_rdData),
    .io_ctrl_rs1En(regs_io_ctrl_rs1En),
    .io_ctrl_rs2En(regs_io_ctrl_rs2En),
    .io_ctrl_rs1Addr(regs_io_ctrl_rs1Addr),
    .io_ctrl_rs2Addr(regs_io_ctrl_rs2Addr),
    .rf_10(regs_rf_10)
  );
  ImmGen imm ( // @[Decode.scala 36:20]
    .io_inst(imm_io_inst),
    .io_immOp(imm_io_immOp),
    .io_imm(imm_io_imm)
  );
  ContrGen con ( // @[Decode.scala 37:20]
    .io_inst(con_io_inst),
    .io_branch(con_io_branch),
    .io_immOp(con_io_immOp),
    .io_rdEn(con_io_rdEn),
    .io_rdAddr(con_io_rdAddr),
    .io_typeL(con_io_typeL),
    .io_aluCtr_aluA(con_io_aluCtr_aluA),
    .io_aluCtr_aluB(con_io_aluCtr_aluB),
    .io_aluCtr_aluOp(con_io_aluCtr_aluOp),
    .io_memCtr_memtoReg(con_io_memCtr_memtoReg),
    .io_memCtr_memWr(con_io_memCtr_memWr),
    .io_memCtr_memOP(con_io_memCtr_memOP),
    .io_regCtrl_rs1En(con_io_regCtrl_rs1En),
    .io_regCtrl_rs2En(con_io_regCtrl_rs2En),
    .io_regCtrl_rs1Addr(con_io_regCtrl_rs1Addr),
    .io_regCtrl_rs2Addr(con_io_regCtrl_rs2Addr)
  );
  assign io_bubbleId = rdRs1HitEx | rdRs2HitEx; // @[Decode.scala 111:30]
  assign io_out_valid = io_in_valid; // @[Decode.scala 90:19]
  assign io_out_pc = io_in_pc; // @[Decode.scala 91:19]
  assign io_out_inst = io_in_inst; // @[Decode.scala 92:19]
  assign io_out_typeL = con_io_typeL; // @[Decode.scala 93:19]
  assign io_out_aluA = con_io_aluCtr_aluA; // @[Decode.scala 94:19]
  assign io_out_aluB = con_io_aluCtr_aluB; // @[Decode.scala 95:19]
  assign io_out_aluOp = con_io_aluCtr_aluOp; // @[Decode.scala 96:19]
  assign io_out_branch = con_io_branch; // @[Decode.scala 97:19]
  assign io_out_memtoReg = con_io_memCtr_memtoReg; // @[Decode.scala 98:19]
  assign io_out_memWr = con_io_memCtr_memWr; // @[Decode.scala 99:19]
  assign io_out_memOp = con_io_memCtr_memOP; // @[Decode.scala 100:19]
  assign io_out_rdEn = con_io_rdEn; // @[Decode.scala 101:19]
  assign io_out_rdAddr = con_io_rdAddr; // @[Decode.scala 102:19]
  assign io_out_rs1Data = con_io_regCtrl_rs1En ? _rs1Data_T_2 : 64'h0; // @[Decode.scala 60:20]
  assign io_out_rs2Data = con_io_regCtrl_rs2En ? _rs2Data_T_2 : 64'h0; // @[Decode.scala 65:20]
  assign io_out_imm = imm_io_imm; // @[Decode.scala 105:19]
  assign rf_10 = regs_rf_10;
  assign regs_clock = clock;
  assign regs_reset = reset;
  assign regs_io_rdEn = io_rdEn; // @[Decode.scala 40:16]
  assign regs_io_rdAddr = {{27'd0}, io_rdAddr}; // @[Decode.scala 41:18]
  assign regs_io_rdData = io_rdData; // @[Decode.scala 42:18]
  assign regs_io_ctrl_rs1En = con_io_regCtrl_rs1En; // @[Decode.scala 39:16]
  assign regs_io_ctrl_rs2En = con_io_regCtrl_rs2En; // @[Decode.scala 39:16]
  assign regs_io_ctrl_rs1Addr = con_io_regCtrl_rs1Addr; // @[Decode.scala 39:16]
  assign regs_io_ctrl_rs2Addr = con_io_regCtrl_rs2Addr; // @[Decode.scala 39:16]
  assign imm_io_inst = io_in_inst; // @[Decode.scala 44:15]
  assign imm_io_immOp = con_io_immOp; // @[Decode.scala 45:16]
  assign con_io_inst = io_in_inst; // @[Decode.scala 46:15]
endmodule
module ALU(
  input  [1:0]  io_memtoReg,
  input  [31:0] io_pc,
  output [63:0] io_aluRes,
  output        io_less,
  output        io_zero,
  input         ctrl_aluA,
  input  [1:0]  ctrl_aluB,
  input  [3:0]  ctrl_aluOp,
  input  [63:0] data_rData1,
  input  [63:0] data_rData2,
  input  [63:0] data_imm
);
  wire [63:0] Asrc = ~ctrl_aluA ? data_rData1 : {{32'd0}, io_pc}; // @[ALU.scala 23:19]
  wire  instW = io_memtoReg[1]; // @[ALU.scala 25:28]
  wire  in1_signBit = Asrc[31]; // @[BitUtils.scala 18:20]
  wire [31:0] _in1_T_3 = in1_signBit ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _in1_T_4 = {_in1_T_3,Asrc[31:0]}; // @[Cat.scala 31:58]
  wire [63:0] _in1_T_6 = {32'h0,Asrc[31:0]}; // @[Cat.scala 31:58]
  wire [63:0] _in1_T_7 = ctrl_aluOp == 4'hd ? _in1_T_4 : _in1_T_6; // @[ALU.scala 26:30]
  wire [63:0] in1 = instW ? _in1_T_7 : Asrc; // @[ALU.scala 26:18]
  wire [63:0] _in2_T_1 = 2'h1 == ctrl_aluB ? data_imm : data_rData2; // @[Mux.scala 81:58]
  wire [63:0] _in2_T_3 = 2'h2 == ctrl_aluB ? 64'h4 : _in2_T_1; // @[Mux.scala 81:58]
  wire [63:0] in2 = 2'h3 == ctrl_aluB ? 64'h0 : _in2_T_3; // @[Mux.scala 81:58]
  wire [5:0] shamt = instW ? {{1'd0}, in2[4:0]} : in2[5:0]; // @[ALU.scala 36:20]
  wire [63:0] addRes = in1 + in2; // @[ALU.scala 38:25]
  wire [63:0] subRes = in1 - in2; // @[ALU.scala 39:25]
  wire [63:0] xorRes = in1 ^ in2; // @[ALU.scala 40:25]
  wire [63:0] orRes = in1 | in2; // @[ALU.scala 41:25]
  wire [63:0] andRes = in1 & in2; // @[ALU.scala 42:25]
  wire [126:0] _GEN_0 = {{63'd0}, in1}; // @[ALU.scala 43:28]
  wire [126:0] _sLRes_T = _GEN_0 << shamt; // @[ALU.scala 43:28]
  wire [63:0] sLRes = _sLRes_T[63:0]; // @[ALU.scala 43:37]
  wire [63:0] sRLRes = in1 >> shamt; // @[ALU.scala 44:27]
  wire [63:0] _sRARes_T = instW ? _in1_T_7 : Asrc; // @[ALU.scala 45:33]
  wire [63:0] sRARes = $signed(_sRARes_T) >>> shamt; // @[ALU.scala 45:52]
  wire [63:0] _sLTRes_T_1 = 2'h3 == ctrl_aluB ? 64'h0 : _in2_T_3; // @[ALU.scala 47:48]
  wire  sLTRes = $signed(_sRARes_T) < $signed(_sLTRes_T_1); // @[ALU.scala 47:36]
  wire  sLTURes = in1 < in2; // @[ALU.scala 48:27]
  wire [63:0] remwRes = $signed(_sRARes_T) % $signed(_sLTRes_T_1); // @[ALU.scala 50:48]
  wire [63:0] divRes = in1 / in2; // @[ALU.scala 51:27]
  wire [127:0] mulRes = in1 * in2; // @[ALU.scala 52:27]
  wire [63:0] _aluResult_T_1 = 4'h0 == ctrl_aluOp ? addRes : 64'h0; // @[Mux.scala 81:58]
  wire [63:0] _aluResult_T_3 = 4'h8 == ctrl_aluOp ? subRes : _aluResult_T_1; // @[Mux.scala 81:58]
  wire [63:0] _aluResult_T_5 = 4'h9 == ctrl_aluOp ? subRes : _aluResult_T_3; // @[Mux.scala 81:58]
  wire [63:0] _aluResult_T_7 = 4'h2 == ctrl_aluOp ? {{63'd0}, sLTRes} : _aluResult_T_5; // @[Mux.scala 81:58]
  wire [63:0] _aluResult_T_9 = 4'ha == ctrl_aluOp ? {{63'd0}, sLTURes} : _aluResult_T_7; // @[Mux.scala 81:58]
  wire [63:0] _aluResult_T_11 = 4'h5 == ctrl_aluOp ? sRLRes : _aluResult_T_9; // @[Mux.scala 81:58]
  wire [63:0] _aluResult_T_13 = 4'hd == ctrl_aluOp ? sRARes : _aluResult_T_11; // @[Mux.scala 81:58]
  wire [63:0] _aluResult_T_15 = 4'h1 == ctrl_aluOp ? sLRes : _aluResult_T_13; // @[Mux.scala 81:58]
  wire [63:0] _aluResult_T_17 = 4'h3 == ctrl_aluOp ? in2 : _aluResult_T_15; // @[Mux.scala 81:58]
  wire [63:0] _aluResult_T_19 = 4'hb == ctrl_aluOp ? remwRes : _aluResult_T_17; // @[Mux.scala 81:58]
  wire [63:0] _aluResult_T_21 = 4'h4 == ctrl_aluOp ? xorRes : _aluResult_T_19; // @[Mux.scala 81:58]
  wire [63:0] _aluResult_T_23 = 4'hc == ctrl_aluOp ? divRes : _aluResult_T_21; // @[Mux.scala 81:58]
  wire [63:0] _aluResult_T_25 = 4'h6 == ctrl_aluOp ? orRes : _aluResult_T_23; // @[Mux.scala 81:58]
  wire [127:0] _aluResult_T_27 = 4'he == ctrl_aluOp ? mulRes : {{64'd0}, _aluResult_T_25}; // @[Mux.scala 81:58]
  wire [127:0] aluResult = 4'h7 == ctrl_aluOp ? {{64'd0}, andRes} : _aluResult_T_27; // @[Mux.scala 81:58]
  wire  io_aluRes_signBit = aluResult[31]; // @[BitUtils.scala 18:20]
  wire [31:0] _io_aluRes_T_2 = io_aluRes_signBit ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _io_aluRes_T_3 = {_io_aluRes_T_2,aluResult[31:0]}; // @[Cat.scala 31:58]
  wire [127:0] _io_aluRes_T_4 = instW ? {{64'd0}, _io_aluRes_T_3} : aluResult; // @[ALU.scala 80:21]
  assign io_aluRes = _io_aluRes_T_4[63:0]; // @[ALU.scala 80:15]
  assign io_less = ctrl_aluOp[3] ? sLTURes : sLTRes; // @[ALU.scala 78:19]
  assign io_zero = aluResult == 128'h0; // @[ALU.scala 79:27]
endmodule
module NextPC(
  input  [31:0] io_pc,
  input  [63:0] io_imm,
  input  [63:0] io_rs1Data,
  input  [2:0]  io_branch,
  input         io_less,
  input         io_zero,
  output [31:0] io_nextPC,
  output [1:0]  io_pcSrc
);
  wire  less = io_branch == 3'h7 ? ~io_less : io_less; // @[NextPC.scala 23:17]
  wire [3:0] _pcSrc_T_1 = {io_branch,io_zero}; // @[NextPC.scala 26:43]
  wire [3:0] _pcSrc_T_7 = {io_branch,less}; // @[NextPC.scala 27:20]
  wire  _pcSrc_T_8 = _pcSrc_T_7 == 4'hc; // @[NextPC.scala 27:28]
  wire  _pcSrc_T_9 = io_branch == 3'h0 | _pcSrc_T_1 == 4'h8 | _pcSrc_T_1 == 4'hb | _pcSrc_T_8; // @[NextPC.scala 26:109]
  wire  _pcSrc_T_12 = _pcSrc_T_9 | _pcSrc_T_7 == 4'he; // @[NextPC.scala 27:43]
  wire  _pcSrc_T_21 = _pcSrc_T_7 == 4'hd; // @[NextPC.scala 29:28]
  wire  _pcSrc_T_22 = io_branch == 3'h1 | _pcSrc_T_1 == 4'h9 | _pcSrc_T_1 == 4'ha | _pcSrc_T_21; // @[NextPC.scala 28:108]
  wire  _pcSrc_T_25 = _pcSrc_T_22 | _pcSrc_T_7 == 4'hf; // @[NextPC.scala 29:43]
  wire  _pcSrc_T_26 = io_branch == 3'h2; // @[NextPC.scala 30:16]
  wire [1:0] _pcSrc_T_27 = _pcSrc_T_26 ? 2'h3 : 2'h1; // @[Mux.scala 101:16]
  wire [1:0] _pcSrc_T_28 = _pcSrc_T_25 ? 2'h2 : _pcSrc_T_27; // @[Mux.scala 101:16]
  wire [1:0] pcSrc = _pcSrc_T_12 ? 2'h0 : _pcSrc_T_28; // @[Mux.scala 101:16]
  wire [31:0] _io_nextPC_T_1 = io_pc + 32'h4; // @[NextPC.scala 34:23]
  wire [63:0] _GEN_0 = {{32'd0}, io_pc}; // @[NextPC.scala 35:23]
  wire [63:0] _io_nextPC_T_3 = _GEN_0 + io_imm; // @[NextPC.scala 35:23]
  wire [63:0] _io_nextPC_T_5 = io_rs1Data + io_imm; // @[NextPC.scala 36:28]
  wire [31:0] _io_nextPC_T_7 = 2'h0 == pcSrc ? _io_nextPC_T_1 : 32'h80000000; // @[Mux.scala 81:58]
  wire [63:0] _io_nextPC_T_9 = 2'h2 == pcSrc ? _io_nextPC_T_3 : {{32'd0}, _io_nextPC_T_7}; // @[Mux.scala 81:58]
  wire [63:0] _io_nextPC_T_11 = 2'h3 == pcSrc ? _io_nextPC_T_5 : _io_nextPC_T_9; // @[Mux.scala 81:58]
  assign io_nextPC = _io_nextPC_T_11[31:0]; // @[NextPC.scala 33:13]
  assign io_pcSrc = _pcSrc_T_12 ? 2'h0 : _pcSrc_T_28; // @[Mux.scala 101:16]
endmodule
module Execution(
  input         io_in_valid,
  input  [31:0] io_in_pc,
  input  [31:0] io_in_inst,
  input         io_in_typeL,
  input         io_in_aluA,
  input  [1:0]  io_in_aluB,
  input  [3:0]  io_in_aluOp,
  input  [2:0]  io_in_branch,
  input  [1:0]  io_in_memtoReg,
  input         io_in_memWr,
  input  [2:0]  io_in_memOp,
  input         io_in_rdEn,
  input  [4:0]  io_in_rdAddr,
  input  [63:0] io_in_rs1Data,
  input  [63:0] io_in_rs2Data,
  input  [63:0] io_in_imm,
  output        io_out_valid,
  output [31:0] io_out_pc,
  output [31:0] io_out_inst,
  output        io_out_typeL,
  output        io_out_aluA,
  output [1:0]  io_out_aluB,
  output [3:0]  io_out_aluOp,
  output [2:0]  io_out_branch,
  output [1:0]  io_out_memtoReg,
  output        io_out_memWr,
  output [2:0]  io_out_memOp,
  output        io_out_rdEn,
  output [4:0]  io_out_rdAddr,
  output [63:0] io_out_rs1Data,
  output [63:0] io_out_rs2Data,
  output [63:0] io_out_imm,
  output [63:0] io_out_aluRes,
  output        io_exeRdEn,
  output [4:0]  io_exeRdAddr,
  output [63:0] io_exeRdData,
  output        io_bubbleEx,
  output [1:0]  io_pcSrc,
  output [31:0] io_nextPC
);
  wire [1:0] alu_io_memtoReg; // @[Execution.scala 20:21]
  wire [31:0] alu_io_pc; // @[Execution.scala 20:21]
  wire [63:0] alu_io_aluRes; // @[Execution.scala 20:21]
  wire  alu_io_less; // @[Execution.scala 20:21]
  wire  alu_io_zero; // @[Execution.scala 20:21]
  wire  alu_ctrl_aluA; // @[Execution.scala 20:21]
  wire [1:0] alu_ctrl_aluB; // @[Execution.scala 20:21]
  wire [3:0] alu_ctrl_aluOp; // @[Execution.scala 20:21]
  wire [63:0] alu_data_rData1; // @[Execution.scala 20:21]
  wire [63:0] alu_data_rData2; // @[Execution.scala 20:21]
  wire [63:0] alu_data_imm; // @[Execution.scala 20:21]
  wire [31:0] nextPC_io_pc; // @[Execution.scala 21:24]
  wire [63:0] nextPC_io_imm; // @[Execution.scala 21:24]
  wire [63:0] nextPC_io_rs1Data; // @[Execution.scala 21:24]
  wire [2:0] nextPC_io_branch; // @[Execution.scala 21:24]
  wire  nextPC_io_less; // @[Execution.scala 21:24]
  wire  nextPC_io_zero; // @[Execution.scala 21:24]
  wire [31:0] nextPC_io_nextPC; // @[Execution.scala 21:24]
  wire [1:0] nextPC_io_pcSrc; // @[Execution.scala 21:24]
  ALU alu ( // @[Execution.scala 20:21]
    .io_memtoReg(alu_io_memtoReg),
    .io_pc(alu_io_pc),
    .io_aluRes(alu_io_aluRes),
    .io_less(alu_io_less),
    .io_zero(alu_io_zero),
    .ctrl_aluA(alu_ctrl_aluA),
    .ctrl_aluB(alu_ctrl_aluB),
    .ctrl_aluOp(alu_ctrl_aluOp),
    .data_rData1(alu_data_rData1),
    .data_rData2(alu_data_rData2),
    .data_imm(alu_data_imm)
  );
  NextPC nextPC ( // @[Execution.scala 21:24]
    .io_pc(nextPC_io_pc),
    .io_imm(nextPC_io_imm),
    .io_rs1Data(nextPC_io_rs1Data),
    .io_branch(nextPC_io_branch),
    .io_less(nextPC_io_less),
    .io_zero(nextPC_io_zero),
    .io_nextPC(nextPC_io_nextPC),
    .io_pcSrc(nextPC_io_pcSrc)
  );
  assign io_out_valid = io_in_valid; // @[Execution.scala 60:19]
  assign io_out_pc = io_in_pc; // @[Execution.scala 61:19]
  assign io_out_inst = io_in_inst; // @[Execution.scala 62:19]
  assign io_out_typeL = io_in_typeL; // @[Execution.scala 63:19]
  assign io_out_aluA = io_in_aluA; // @[Execution.scala 64:19]
  assign io_out_aluB = io_in_aluB; // @[Execution.scala 65:19]
  assign io_out_aluOp = io_in_aluOp; // @[Execution.scala 66:19]
  assign io_out_branch = io_in_branch; // @[Execution.scala 67:19]
  assign io_out_memtoReg = io_in_memtoReg; // @[Execution.scala 68:19]
  assign io_out_memWr = io_in_memWr; // @[Execution.scala 69:19]
  assign io_out_memOp = io_in_memOp; // @[Execution.scala 70:19]
  assign io_out_rdEn = io_in_rdEn; // @[Execution.scala 71:19]
  assign io_out_rdAddr = io_in_rdAddr; // @[Execution.scala 72:19]
  assign io_out_rs1Data = io_in_rs1Data; // @[Execution.scala 73:19]
  assign io_out_rs2Data = io_in_rs2Data; // @[Execution.scala 74:19]
  assign io_out_imm = io_in_imm; // @[Execution.scala 75:19]
  assign io_out_aluRes = alu_io_aluRes; // @[Execution.scala 78:19]
  assign io_exeRdEn = io_in_rdEn; // @[Execution.scala 81:14]
  assign io_exeRdAddr = io_in_rdAddr; // @[Execution.scala 82:16]
  assign io_exeRdData = alu_io_aluRes; // @[Execution.scala 83:16]
  assign io_bubbleEx = io_in_typeL; // @[Execution.scala 85:15]
  assign io_pcSrc = nextPC_io_pcSrc; // @[Execution.scala 87:12]
  assign io_nextPC = nextPC_io_nextPC; // @[Execution.scala 88:13]
  assign alu_io_memtoReg = io_in_memtoReg; // @[Execution.scala 28:21]
  assign alu_io_pc = io_in_pc; // @[Execution.scala 29:15]
  assign alu_ctrl_aluA = io_in_aluA; // @[Execution.scala 22:25]
  assign alu_ctrl_aluB = io_in_aluB; // @[Execution.scala 23:25]
  assign alu_ctrl_aluOp = io_in_aluOp; // @[Execution.scala 24:26]
  assign alu_data_rData1 = io_in_rs1Data; // @[Execution.scala 25:27]
  assign alu_data_rData2 = io_in_rs2Data; // @[Execution.scala 26:27]
  assign alu_data_imm = io_in_imm; // @[Execution.scala 27:24]
  assign nextPC_io_pc = io_in_pc; // @[Execution.scala 31:18]
  assign nextPC_io_imm = io_in_imm; // @[Execution.scala 32:19]
  assign nextPC_io_rs1Data = io_in_rs1Data; // @[Execution.scala 33:23]
  assign nextPC_io_branch = io_in_branch; // @[Execution.scala 34:22]
  assign nextPC_io_less = alu_io_less; // @[Execution.scala 35:20]
  assign nextPC_io_zero = alu_io_zero; // @[Execution.scala 36:20]
endmodule
module DataMem(
  input          clock,
  input          reset,
  output         io_dmem_data_valid,
  input          io_dmem_data_ready,
  output         io_dmem_data_req,
  output [31:0]  io_dmem_data_addr,
  output [1:0]   io_dmem_data_size,
  output [7:0]   io_dmem_data_strb,
  input  [63:0]  io_dmem_data_read,
  output [127:0] io_dmem_data_write,
  input          io_in_valid,
  input  [31:0]  io_in_pc,
  input  [31:0]  io_in_inst,
  input          io_in_typeL,
  input          io_in_aluA,
  input  [1:0]   io_in_aluB,
  input  [3:0]   io_in_aluOp,
  input  [2:0]   io_in_branch,
  input  [1:0]   io_in_memtoReg,
  input          io_in_memWr,
  input  [2:0]   io_in_memOp,
  input          io_in_rdEn,
  input  [4:0]   io_in_rdAddr,
  input  [63:0]  io_in_rs1Data,
  input  [63:0]  io_in_rs2Data,
  input  [63:0]  io_in_imm,
  input  [63:0]  io_in_aluRes,
  output         io_out_valid,
  output [31:0]  io_out_pc,
  output [31:0]  io_out_inst,
  output         io_out_typeL,
  output         io_out_aluA,
  output [1:0]   io_out_aluB,
  output [3:0]   io_out_aluOp,
  output [2:0]   io_out_branch,
  output [1:0]   io_out_memtoReg,
  output         io_out_memWr,
  output [2:0]   io_out_memOp,
  output         io_out_rdEn,
  output [4:0]   io_out_rdAddr,
  output [63:0]  io_out_rs1Data,
  output [63:0]  io_out_rs2Data,
  output [63:0]  io_out_imm,
  output [63:0]  io_out_aluRes,
  output [63:0]  io_out_memData,
  input          io_IFReady,
  output         io_memRdEn,
  output [4:0]   io_memRdAddr,
  output [63:0]  io_memRdData,
  output         io_memDone
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  _dmemEn_T_6 = io_in_memtoReg == 2'h1 | io_in_memWr; // @[DataMem.scala 39:43]
  wire  dmemEn = ~(io_in_aluRes < 64'h80000000 | io_in_aluRes > 64'h88000000) & _dmemEn_T_6; // @[DataMem.scala 38:72]
  reg  dmemDone; // @[DataMem.scala 43:25]
  reg [31:0] inst; // @[DataMem.scala 44:17]
  wire  _GEN_0 = inst != io_in_inst ? 1'h0 : dmemDone; // @[DataMem.scala 49:37 50:14 43:25]
  wire  _GEN_1 = io_dmem_data_ready | _GEN_0; // @[DataMem.scala 47:29 48:14]
  wire  dmemFire = io_dmem_data_valid & io_dmem_data_ready; // @[DataMem.scala 55:37]
  wire [63:0] _GEN_3 = io_in_aluRes % 64'h10; // @[DataMem.scala 56:27]
  wire [4:0] alignBits = _GEN_3[4:0]; // @[DataMem.scala 56:27]
  wire [8:0] _io_dmem_data_write_T = alignBits * 4'h8; // @[DataMem.scala 58:48]
  wire [574:0] _GEN_4 = {{511'd0}, io_in_rs2Data}; // @[DataMem.scala 58:35]
  wire [574:0] _io_dmem_data_write_T_1 = _GEN_4 << _io_dmem_data_write_T; // @[DataMem.scala 58:35]
  wire [1:0] _io_dmem_data_strb_T_1 = 5'h1 == alignBits ? 2'h2 : 2'h1; // @[Mux.scala 81:58]
  wire [2:0] _io_dmem_data_strb_T_3 = 5'h2 == alignBits ? 3'h4 : {{1'd0}, _io_dmem_data_strb_T_1}; // @[Mux.scala 81:58]
  wire [3:0] _io_dmem_data_strb_T_5 = 5'h3 == alignBits ? 4'h8 : {{1'd0}, _io_dmem_data_strb_T_3}; // @[Mux.scala 81:58]
  wire [4:0] _io_dmem_data_strb_T_7 = 5'h4 == alignBits ? 5'h10 : {{1'd0}, _io_dmem_data_strb_T_5}; // @[Mux.scala 81:58]
  wire [5:0] _io_dmem_data_strb_T_9 = 5'h5 == alignBits ? 6'h20 : {{1'd0}, _io_dmem_data_strb_T_7}; // @[Mux.scala 81:58]
  wire [6:0] _io_dmem_data_strb_T_11 = 5'h6 == alignBits ? 7'h40 : {{1'd0}, _io_dmem_data_strb_T_9}; // @[Mux.scala 81:58]
  wire [7:0] _io_dmem_data_strb_T_13 = 5'h7 == alignBits ? 8'h80 : {{1'd0}, _io_dmem_data_strb_T_11}; // @[Mux.scala 81:58]
  wire [7:0] _io_dmem_data_strb_T_15 = 5'h9 == alignBits ? 8'h2 : _io_dmem_data_strb_T_13; // @[Mux.scala 81:58]
  wire [7:0] _io_dmem_data_strb_T_17 = 5'ha == alignBits ? 8'h4 : _io_dmem_data_strb_T_15; // @[Mux.scala 81:58]
  wire [7:0] _io_dmem_data_strb_T_19 = 5'hb == alignBits ? 8'h8 : _io_dmem_data_strb_T_17; // @[Mux.scala 81:58]
  wire [7:0] _io_dmem_data_strb_T_21 = 5'hc == alignBits ? 8'h10 : _io_dmem_data_strb_T_19; // @[Mux.scala 81:58]
  wire [7:0] _io_dmem_data_strb_T_23 = 5'hd == alignBits ? 8'h20 : _io_dmem_data_strb_T_21; // @[Mux.scala 81:58]
  wire [7:0] _io_dmem_data_strb_T_25 = 5'he == alignBits ? 8'h40 : _io_dmem_data_strb_T_23; // @[Mux.scala 81:58]
  wire [7:0] _io_dmem_data_strb_T_27 = 5'hf == alignBits ? 8'h80 : _io_dmem_data_strb_T_25; // @[Mux.scala 81:58]
  wire [3:0] _io_dmem_data_strb_T_29 = 5'h2 == alignBits ? 4'hc : 4'h3; // @[Mux.scala 81:58]
  wire [5:0] _io_dmem_data_strb_T_31 = 5'h4 == alignBits ? 6'h30 : {{2'd0}, _io_dmem_data_strb_T_29}; // @[Mux.scala 81:58]
  wire [7:0] _io_dmem_data_strb_T_33 = 5'h6 == alignBits ? 8'hc0 : {{2'd0}, _io_dmem_data_strb_T_31}; // @[Mux.scala 81:58]
  wire [7:0] _io_dmem_data_strb_T_35 = 5'ha == alignBits ? 8'hc : _io_dmem_data_strb_T_33; // @[Mux.scala 81:58]
  wire [7:0] _io_dmem_data_strb_T_37 = 5'hc == alignBits ? 8'h30 : _io_dmem_data_strb_T_35; // @[Mux.scala 81:58]
  wire [7:0] _io_dmem_data_strb_T_39 = 5'he == alignBits ? 8'hc0 : _io_dmem_data_strb_T_37; // @[Mux.scala 81:58]
  wire [7:0] _io_dmem_data_strb_T_43 = alignBits == 5'h0 | alignBits == 5'h8 ? 8'hf : 8'hf0; // @[DataMem.scala 88:22]
  wire [7:0] _io_dmem_data_strb_T_45 = 3'h0 == io_in_memOp ? _io_dmem_data_strb_T_27 : 8'h0; // @[Mux.scala 81:58]
  wire [7:0] _io_dmem_data_strb_T_47 = 3'h1 == io_in_memOp ? _io_dmem_data_strb_T_39 : _io_dmem_data_strb_T_45; // @[Mux.scala 81:58]
  wire [7:0] _io_dmem_data_strb_T_49 = 3'h2 == io_in_memOp ? _io_dmem_data_strb_T_43 : _io_dmem_data_strb_T_47; // @[Mux.scala 81:58]
  wire [7:0] _io_dmem_data_strb_T_51 = 3'h3 == io_in_memOp ? 8'hff : _io_dmem_data_strb_T_49; // @[Mux.scala 81:58]
  reg [63:0] rdata; // @[DataMem.scala 93:22]
  wire  memAxi = dmemEn & ~dmemFire; // @[DataMem.scala 98:27]
  wire  rData_signBit = rdata[7]; // @[BitUtils.scala 18:20]
  wire [55:0] _rData_T_2 = rData_signBit ? 56'hffffffffffffff : 56'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _rData_T_3 = {_rData_T_2,rdata[7:0]}; // @[Cat.scala 31:58]
  wire  rData_signBit_1 = rdata[15]; // @[BitUtils.scala 18:20]
  wire [47:0] _rData_T_6 = rData_signBit_1 ? 48'hffffffffffff : 48'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _rData_T_7 = {_rData_T_6,rdata[15:0]}; // @[Cat.scala 31:58]
  wire  rData_signBit_2 = rdata[31]; // @[BitUtils.scala 18:20]
  wire [31:0] _rData_T_10 = rData_signBit_2 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _rData_T_11 = {_rData_T_10,rdata[31:0]}; // @[Cat.scala 31:58]
  wire [63:0] _rData_T_13 = {56'h0,rdata[7:0]}; // @[Cat.scala 31:58]
  wire [63:0] _rData_T_15 = {48'h0,rdata[15:0]}; // @[Cat.scala 31:58]
  wire [63:0] _rData_T_17 = {32'h0,rdata[31:0]}; // @[Cat.scala 31:58]
  wire [63:0] _rData_T_19 = 3'h0 == io_in_memOp ? _rData_T_3 : 64'h0; // @[Mux.scala 81:58]
  wire [63:0] _rData_T_21 = 3'h1 == io_in_memOp ? _rData_T_7 : _rData_T_19; // @[Mux.scala 81:58]
  wire [63:0] _rData_T_23 = 3'h2 == io_in_memOp ? _rData_T_11 : _rData_T_21; // @[Mux.scala 81:58]
  wire [63:0] _rData_T_25 = 3'h3 == io_in_memOp ? rdata : _rData_T_23; // @[Mux.scala 81:58]
  wire [63:0] _rData_T_27 = 3'h4 == io_in_memOp ? _rData_T_13 : _rData_T_25; // @[Mux.scala 81:58]
  wire [63:0] _rData_T_29 = 3'h5 == io_in_memOp ? _rData_T_15 : _rData_T_27; // @[Mux.scala 81:58]
  wire [63:0] rData = 3'h6 == io_in_memOp ? _rData_T_17 : _rData_T_29; // @[Mux.scala 81:58]
  wire  _data_size_T_7 = 3'h5 == io_in_memOp | 3'h1 == io_in_memOp; // @[Mux.scala 81:58]
  wire [1:0] _data_size_T_9 = 3'h3 == io_in_memOp ? 2'h3 : {{1'd0}, _data_size_T_7}; // @[Mux.scala 81:58]
  wire [1:0] _data_size_T_11 = 3'h2 == io_in_memOp ? 2'h2 : _data_size_T_9; // @[Mux.scala 81:58]
  wire [63:0] memData = io_in_memWr ? 64'h0 : rData; // @[DataMem.scala 155:18]
  wire  resW_signBit = io_in_aluRes[31]; // @[BitUtils.scala 18:20]
  wire [31:0] _resW_T_2 = resW_signBit ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] resW = {_resW_T_2,io_in_aluRes[31:0]}; // @[Cat.scala 31:58]
  wire [63:0] _memBPData_T_1 = 2'h0 == io_in_memtoReg ? io_in_aluRes : 64'h0; // @[Mux.scala 81:58]
  wire [63:0] _memBPData_T_3 = 2'h1 == io_in_memtoReg ? memData : _memBPData_T_1; // @[Mux.scala 81:58]
  assign io_dmem_data_valid = dmemEn & ~io_IFReady & ~dmemDone; // @[DataMem.scala 53:47]
  assign io_dmem_data_req = io_in_memWr; // @[DataMem.scala 59:26]
  assign io_dmem_data_addr = io_in_aluRes[31:0]; // @[DataMem.scala 41:21]
  assign io_dmem_data_size = 3'h6 == io_in_memOp ? 2'h2 : _data_size_T_11; // @[Mux.scala 81:58]
  assign io_dmem_data_strb = io_in_typeL ? 8'h0 : _io_dmem_data_strb_T_51; // @[DataMem.scala 61:27]
  assign io_dmem_data_write = _io_dmem_data_write_T_1[127:0]; // @[DataMem.scala 58:22]
  assign io_out_valid = io_in_valid; // @[DataMem.scala 186:19]
  assign io_out_pc = io_in_pc; // @[DataMem.scala 187:19]
  assign io_out_inst = io_in_inst; // @[DataMem.scala 188:19]
  assign io_out_typeL = io_in_typeL; // @[DataMem.scala 189:19]
  assign io_out_aluA = io_in_aluA; // @[DataMem.scala 190:19]
  assign io_out_aluB = io_in_aluB; // @[DataMem.scala 191:19]
  assign io_out_aluOp = io_in_aluOp; // @[DataMem.scala 192:19]
  assign io_out_branch = io_in_branch; // @[DataMem.scala 193:19]
  assign io_out_memtoReg = io_in_memtoReg; // @[DataMem.scala 194:19]
  assign io_out_memWr = io_in_memWr; // @[DataMem.scala 195:19]
  assign io_out_memOp = io_in_memOp; // @[DataMem.scala 196:19]
  assign io_out_rdEn = io_in_rdEn; // @[DataMem.scala 197:19]
  assign io_out_rdAddr = io_in_rdAddr; // @[DataMem.scala 198:19]
  assign io_out_rs1Data = io_in_rs1Data; // @[DataMem.scala 199:19]
  assign io_out_rs2Data = io_in_rs2Data; // @[DataMem.scala 200:19]
  assign io_out_imm = io_in_imm; // @[DataMem.scala 201:19]
  assign io_out_aluRes = io_in_aluRes; // @[DataMem.scala 204:19]
  assign io_out_memData = io_in_memWr ? 64'h0 : rData; // @[DataMem.scala 155:18]
  assign io_memRdEn = io_in_rdEn; // @[DataMem.scala 207:14]
  assign io_memRdAddr = io_in_rdAddr; // @[DataMem.scala 208:16]
  assign io_memRdData = 2'h2 == io_in_memtoReg ? resW : _memBPData_T_3; // @[Mux.scala 81:58]
  assign io_memDone = ~io_in_typeL ? ~memAxi | io_IFReady : dmemDone; // @[DataMem.scala 100:20]
  always @(posedge clock) begin
    if (reset) begin // @[DataMem.scala 43:25]
      dmemDone <= 1'h0; // @[DataMem.scala 43:25]
    end else begin
      dmemDone <= _GEN_1;
    end
    inst <= io_in_inst; // @[DataMem.scala 46:8]
    if (reset) begin // @[DataMem.scala 93:22]
      rdata <= 64'h0; // @[DataMem.scala 93:22]
    end else if (dmemFire) begin // @[DataMem.scala 94:18]
      rdata <= io_dmem_data_read; // @[DataMem.scala 95:11]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  dmemDone = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  inst = _RAND_1[31:0];
  _RAND_2 = {2{`RANDOM}};
  rdata = _RAND_2[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module WriteBack(
  input         io_in_valid,
  input  [31:0] io_in_pc,
  input  [31:0] io_in_inst,
  input  [1:0]  io_in_memtoReg,
  input         io_in_rdEn,
  input  [4:0]  io_in_rdAddr,
  input  [63:0] io_in_aluRes,
  input  [63:0] io_in_memData,
  output [31:0] io_pc,
  output [31:0] io_inst,
  output        io_rdEn,
  output [4:0]  io_rdAddr,
  output [63:0] io_rdData,
  output        io_wbRdEn,
  output [4:0]  io_wbRdAddr,
  output [63:0] io_wbRdData,
  output        io_ready_cmt
);
  wire  resW_signBit = io_in_aluRes[31]; // @[BitUtils.scala 18:20]
  wire [31:0] _resW_T_2 = resW_signBit ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] resW = {_resW_T_2,io_in_aluRes[31:0]}; // @[Cat.scala 31:58]
  wire [63:0] _rdData_T_1 = 2'h0 == io_in_memtoReg ? io_in_aluRes : 64'h0; // @[Mux.scala 81:58]
  wire [63:0] _rdData_T_3 = 2'h1 == io_in_memtoReg ? io_in_memData : _rdData_T_1; // @[Mux.scala 81:58]
  assign io_pc = io_in_pc; // @[WriteBack.scala 32:9]
  assign io_inst = io_in_inst; // @[WriteBack.scala 33:11]
  assign io_rdEn = io_in_rdEn; // @[WriteBack.scala 35:11]
  assign io_rdAddr = io_in_rdAddr; // @[WriteBack.scala 36:13]
  assign io_rdData = 2'h2 == io_in_memtoReg ? resW : _rdData_T_3; // @[Mux.scala 81:58]
  assign io_wbRdEn = io_in_rdEn; // @[WriteBack.scala 40:13]
  assign io_wbRdAddr = io_in_rdAddr; // @[WriteBack.scala 41:15]
  assign io_wbRdData = 2'h2 == io_in_memtoReg ? resW : _rdData_T_3; // @[Mux.scala 81:58]
  assign io_ready_cmt = io_in_inst != 32'h0 & io_in_valid; // @[WriteBack.scala 38:38]
endmodule
module Core(
  input          clock,
  input          reset,
  output         io_imem_inst_valid,
  input          io_imem_inst_ready,
  output [31:0]  io_imem_inst_addr,
  input  [31:0]  io_imem_inst_read,
  output         io_dmem_data_valid,
  input          io_dmem_data_ready,
  output         io_dmem_data_req,
  output [31:0]  io_dmem_data_addr,
  output [1:0]   io_dmem_data_size,
  output [7:0]   io_dmem_data_strb,
  input  [63:0]  io_dmem_data_read,
  output [127:0] io_dmem_data_write
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  wire  IF_clock; // @[Core.scala 14:18]
  wire  IF_reset; // @[Core.scala 14:18]
  wire  IF_io_imem_inst_valid; // @[Core.scala 14:18]
  wire  IF_io_imem_inst_ready; // @[Core.scala 14:18]
  wire [31:0] IF_io_imem_inst_addr; // @[Core.scala 14:18]
  wire [31:0] IF_io_imem_inst_read; // @[Core.scala 14:18]
  wire [1:0] IF_io_pcSrc; // @[Core.scala 14:18]
  wire [31:0] IF_io_nextPC; // @[Core.scala 14:18]
  wire  IF_io_stall; // @[Core.scala 14:18]
  wire  IF_io_memDone; // @[Core.scala 14:18]
  wire  IF_io_out_valid; // @[Core.scala 14:18]
  wire [31:0] IF_io_out_pc; // @[Core.scala 14:18]
  wire [31:0] IF_io_out_inst; // @[Core.scala 14:18]
  wire  IF_io_IFDone; // @[Core.scala 14:18]
  wire  IfRegId_clock; // @[Core.scala 15:23]
  wire  IfRegId_reset; // @[Core.scala 15:23]
  wire  IfRegId_io_in_valid; // @[Core.scala 15:23]
  wire [31:0] IfRegId_io_in_pc; // @[Core.scala 15:23]
  wire [31:0] IfRegId_io_in_inst; // @[Core.scala 15:23]
  wire  IfRegId_io_in_typeL; // @[Core.scala 15:23]
  wire  IfRegId_io_in_aluA; // @[Core.scala 15:23]
  wire [1:0] IfRegId_io_in_aluB; // @[Core.scala 15:23]
  wire [3:0] IfRegId_io_in_aluOp; // @[Core.scala 15:23]
  wire [2:0] IfRegId_io_in_branch; // @[Core.scala 15:23]
  wire [1:0] IfRegId_io_in_memtoReg; // @[Core.scala 15:23]
  wire  IfRegId_io_in_memWr; // @[Core.scala 15:23]
  wire [2:0] IfRegId_io_in_memOp; // @[Core.scala 15:23]
  wire  IfRegId_io_in_rdEn; // @[Core.scala 15:23]
  wire [4:0] IfRegId_io_in_rdAddr; // @[Core.scala 15:23]
  wire [63:0] IfRegId_io_in_rs1Data; // @[Core.scala 15:23]
  wire [63:0] IfRegId_io_in_rs2Data; // @[Core.scala 15:23]
  wire [63:0] IfRegId_io_in_imm; // @[Core.scala 15:23]
  wire [63:0] IfRegId_io_in_aluRes; // @[Core.scala 15:23]
  wire [63:0] IfRegId_io_in_memData; // @[Core.scala 15:23]
  wire  IfRegId_io_out_valid; // @[Core.scala 15:23]
  wire [31:0] IfRegId_io_out_pc; // @[Core.scala 15:23]
  wire [31:0] IfRegId_io_out_inst; // @[Core.scala 15:23]
  wire  IfRegId_io_out_typeL; // @[Core.scala 15:23]
  wire  IfRegId_io_out_aluA; // @[Core.scala 15:23]
  wire [1:0] IfRegId_io_out_aluB; // @[Core.scala 15:23]
  wire [3:0] IfRegId_io_out_aluOp; // @[Core.scala 15:23]
  wire [2:0] IfRegId_io_out_branch; // @[Core.scala 15:23]
  wire [1:0] IfRegId_io_out_memtoReg; // @[Core.scala 15:23]
  wire  IfRegId_io_out_memWr; // @[Core.scala 15:23]
  wire [2:0] IfRegId_io_out_memOp; // @[Core.scala 15:23]
  wire  IfRegId_io_out_rdEn; // @[Core.scala 15:23]
  wire [4:0] IfRegId_io_out_rdAddr; // @[Core.scala 15:23]
  wire [63:0] IfRegId_io_out_rs1Data; // @[Core.scala 15:23]
  wire [63:0] IfRegId_io_out_rs2Data; // @[Core.scala 15:23]
  wire [63:0] IfRegId_io_out_imm; // @[Core.scala 15:23]
  wire [63:0] IfRegId_io_out_aluRes; // @[Core.scala 15:23]
  wire [63:0] IfRegId_io_out_memData; // @[Core.scala 15:23]
  wire  IfRegId_io_flush; // @[Core.scala 15:23]
  wire  IfRegId_io_stall; // @[Core.scala 15:23]
  wire  ID_clock; // @[Core.scala 16:18]
  wire  ID_reset; // @[Core.scala 16:18]
  wire  ID_io_rdEn; // @[Core.scala 16:18]
  wire [4:0] ID_io_rdAddr; // @[Core.scala 16:18]
  wire [63:0] ID_io_rdData; // @[Core.scala 16:18]
  wire  ID_io_in_valid; // @[Core.scala 16:18]
  wire [31:0] ID_io_in_pc; // @[Core.scala 16:18]
  wire [31:0] ID_io_in_inst; // @[Core.scala 16:18]
  wire  ID_io_exeRdEn; // @[Core.scala 16:18]
  wire [4:0] ID_io_exeRdAddr; // @[Core.scala 16:18]
  wire [63:0] ID_io_exeRdData; // @[Core.scala 16:18]
  wire  ID_io_memRdEn; // @[Core.scala 16:18]
  wire [4:0] ID_io_memRdAddr; // @[Core.scala 16:18]
  wire [63:0] ID_io_memRdData; // @[Core.scala 16:18]
  wire  ID_io_wbRdEn; // @[Core.scala 16:18]
  wire [4:0] ID_io_wbRdAddr; // @[Core.scala 16:18]
  wire [63:0] ID_io_wbRdData; // @[Core.scala 16:18]
  wire  ID_io_bubbleId; // @[Core.scala 16:18]
  wire  ID_io_out_valid; // @[Core.scala 16:18]
  wire [31:0] ID_io_out_pc; // @[Core.scala 16:18]
  wire [31:0] ID_io_out_inst; // @[Core.scala 16:18]
  wire  ID_io_out_typeL; // @[Core.scala 16:18]
  wire  ID_io_out_aluA; // @[Core.scala 16:18]
  wire [1:0] ID_io_out_aluB; // @[Core.scala 16:18]
  wire [3:0] ID_io_out_aluOp; // @[Core.scala 16:18]
  wire [2:0] ID_io_out_branch; // @[Core.scala 16:18]
  wire [1:0] ID_io_out_memtoReg; // @[Core.scala 16:18]
  wire  ID_io_out_memWr; // @[Core.scala 16:18]
  wire [2:0] ID_io_out_memOp; // @[Core.scala 16:18]
  wire  ID_io_out_rdEn; // @[Core.scala 16:18]
  wire [4:0] ID_io_out_rdAddr; // @[Core.scala 16:18]
  wire [63:0] ID_io_out_rs1Data; // @[Core.scala 16:18]
  wire [63:0] ID_io_out_rs2Data; // @[Core.scala 16:18]
  wire [63:0] ID_io_out_imm; // @[Core.scala 16:18]
  wire [63:0] ID_rf_10; // @[Core.scala 16:18]
  wire  IdRegEx_clock; // @[Core.scala 17:23]
  wire  IdRegEx_reset; // @[Core.scala 17:23]
  wire  IdRegEx_io_in_valid; // @[Core.scala 17:23]
  wire [31:0] IdRegEx_io_in_pc; // @[Core.scala 17:23]
  wire [31:0] IdRegEx_io_in_inst; // @[Core.scala 17:23]
  wire  IdRegEx_io_in_typeL; // @[Core.scala 17:23]
  wire  IdRegEx_io_in_aluA; // @[Core.scala 17:23]
  wire [1:0] IdRegEx_io_in_aluB; // @[Core.scala 17:23]
  wire [3:0] IdRegEx_io_in_aluOp; // @[Core.scala 17:23]
  wire [2:0] IdRegEx_io_in_branch; // @[Core.scala 17:23]
  wire [1:0] IdRegEx_io_in_memtoReg; // @[Core.scala 17:23]
  wire  IdRegEx_io_in_memWr; // @[Core.scala 17:23]
  wire [2:0] IdRegEx_io_in_memOp; // @[Core.scala 17:23]
  wire  IdRegEx_io_in_rdEn; // @[Core.scala 17:23]
  wire [4:0] IdRegEx_io_in_rdAddr; // @[Core.scala 17:23]
  wire [63:0] IdRegEx_io_in_rs1Data; // @[Core.scala 17:23]
  wire [63:0] IdRegEx_io_in_rs2Data; // @[Core.scala 17:23]
  wire [63:0] IdRegEx_io_in_imm; // @[Core.scala 17:23]
  wire [63:0] IdRegEx_io_in_aluRes; // @[Core.scala 17:23]
  wire [63:0] IdRegEx_io_in_memData; // @[Core.scala 17:23]
  wire  IdRegEx_io_out_valid; // @[Core.scala 17:23]
  wire [31:0] IdRegEx_io_out_pc; // @[Core.scala 17:23]
  wire [31:0] IdRegEx_io_out_inst; // @[Core.scala 17:23]
  wire  IdRegEx_io_out_typeL; // @[Core.scala 17:23]
  wire  IdRegEx_io_out_aluA; // @[Core.scala 17:23]
  wire [1:0] IdRegEx_io_out_aluB; // @[Core.scala 17:23]
  wire [3:0] IdRegEx_io_out_aluOp; // @[Core.scala 17:23]
  wire [2:0] IdRegEx_io_out_branch; // @[Core.scala 17:23]
  wire [1:0] IdRegEx_io_out_memtoReg; // @[Core.scala 17:23]
  wire  IdRegEx_io_out_memWr; // @[Core.scala 17:23]
  wire [2:0] IdRegEx_io_out_memOp; // @[Core.scala 17:23]
  wire  IdRegEx_io_out_rdEn; // @[Core.scala 17:23]
  wire [4:0] IdRegEx_io_out_rdAddr; // @[Core.scala 17:23]
  wire [63:0] IdRegEx_io_out_rs1Data; // @[Core.scala 17:23]
  wire [63:0] IdRegEx_io_out_rs2Data; // @[Core.scala 17:23]
  wire [63:0] IdRegEx_io_out_imm; // @[Core.scala 17:23]
  wire [63:0] IdRegEx_io_out_aluRes; // @[Core.scala 17:23]
  wire [63:0] IdRegEx_io_out_memData; // @[Core.scala 17:23]
  wire  IdRegEx_io_flush; // @[Core.scala 17:23]
  wire  IdRegEx_io_stall; // @[Core.scala 17:23]
  wire  EX_io_in_valid; // @[Core.scala 18:18]
  wire [31:0] EX_io_in_pc; // @[Core.scala 18:18]
  wire [31:0] EX_io_in_inst; // @[Core.scala 18:18]
  wire  EX_io_in_typeL; // @[Core.scala 18:18]
  wire  EX_io_in_aluA; // @[Core.scala 18:18]
  wire [1:0] EX_io_in_aluB; // @[Core.scala 18:18]
  wire [3:0] EX_io_in_aluOp; // @[Core.scala 18:18]
  wire [2:0] EX_io_in_branch; // @[Core.scala 18:18]
  wire [1:0] EX_io_in_memtoReg; // @[Core.scala 18:18]
  wire  EX_io_in_memWr; // @[Core.scala 18:18]
  wire [2:0] EX_io_in_memOp; // @[Core.scala 18:18]
  wire  EX_io_in_rdEn; // @[Core.scala 18:18]
  wire [4:0] EX_io_in_rdAddr; // @[Core.scala 18:18]
  wire [63:0] EX_io_in_rs1Data; // @[Core.scala 18:18]
  wire [63:0] EX_io_in_rs2Data; // @[Core.scala 18:18]
  wire [63:0] EX_io_in_imm; // @[Core.scala 18:18]
  wire  EX_io_out_valid; // @[Core.scala 18:18]
  wire [31:0] EX_io_out_pc; // @[Core.scala 18:18]
  wire [31:0] EX_io_out_inst; // @[Core.scala 18:18]
  wire  EX_io_out_typeL; // @[Core.scala 18:18]
  wire  EX_io_out_aluA; // @[Core.scala 18:18]
  wire [1:0] EX_io_out_aluB; // @[Core.scala 18:18]
  wire [3:0] EX_io_out_aluOp; // @[Core.scala 18:18]
  wire [2:0] EX_io_out_branch; // @[Core.scala 18:18]
  wire [1:0] EX_io_out_memtoReg; // @[Core.scala 18:18]
  wire  EX_io_out_memWr; // @[Core.scala 18:18]
  wire [2:0] EX_io_out_memOp; // @[Core.scala 18:18]
  wire  EX_io_out_rdEn; // @[Core.scala 18:18]
  wire [4:0] EX_io_out_rdAddr; // @[Core.scala 18:18]
  wire [63:0] EX_io_out_rs1Data; // @[Core.scala 18:18]
  wire [63:0] EX_io_out_rs2Data; // @[Core.scala 18:18]
  wire [63:0] EX_io_out_imm; // @[Core.scala 18:18]
  wire [63:0] EX_io_out_aluRes; // @[Core.scala 18:18]
  wire  EX_io_exeRdEn; // @[Core.scala 18:18]
  wire [4:0] EX_io_exeRdAddr; // @[Core.scala 18:18]
  wire [63:0] EX_io_exeRdData; // @[Core.scala 18:18]
  wire  EX_io_bubbleEx; // @[Core.scala 18:18]
  wire [1:0] EX_io_pcSrc; // @[Core.scala 18:18]
  wire [31:0] EX_io_nextPC; // @[Core.scala 18:18]
  wire  ExRegMem_clock; // @[Core.scala 19:24]
  wire  ExRegMem_reset; // @[Core.scala 19:24]
  wire  ExRegMem_io_in_valid; // @[Core.scala 19:24]
  wire [31:0] ExRegMem_io_in_pc; // @[Core.scala 19:24]
  wire [31:0] ExRegMem_io_in_inst; // @[Core.scala 19:24]
  wire  ExRegMem_io_in_typeL; // @[Core.scala 19:24]
  wire  ExRegMem_io_in_aluA; // @[Core.scala 19:24]
  wire [1:0] ExRegMem_io_in_aluB; // @[Core.scala 19:24]
  wire [3:0] ExRegMem_io_in_aluOp; // @[Core.scala 19:24]
  wire [2:0] ExRegMem_io_in_branch; // @[Core.scala 19:24]
  wire [1:0] ExRegMem_io_in_memtoReg; // @[Core.scala 19:24]
  wire  ExRegMem_io_in_memWr; // @[Core.scala 19:24]
  wire [2:0] ExRegMem_io_in_memOp; // @[Core.scala 19:24]
  wire  ExRegMem_io_in_rdEn; // @[Core.scala 19:24]
  wire [4:0] ExRegMem_io_in_rdAddr; // @[Core.scala 19:24]
  wire [63:0] ExRegMem_io_in_rs1Data; // @[Core.scala 19:24]
  wire [63:0] ExRegMem_io_in_rs2Data; // @[Core.scala 19:24]
  wire [63:0] ExRegMem_io_in_imm; // @[Core.scala 19:24]
  wire [63:0] ExRegMem_io_in_aluRes; // @[Core.scala 19:24]
  wire [63:0] ExRegMem_io_in_memData; // @[Core.scala 19:24]
  wire  ExRegMem_io_out_valid; // @[Core.scala 19:24]
  wire [31:0] ExRegMem_io_out_pc; // @[Core.scala 19:24]
  wire [31:0] ExRegMem_io_out_inst; // @[Core.scala 19:24]
  wire  ExRegMem_io_out_typeL; // @[Core.scala 19:24]
  wire  ExRegMem_io_out_aluA; // @[Core.scala 19:24]
  wire [1:0] ExRegMem_io_out_aluB; // @[Core.scala 19:24]
  wire [3:0] ExRegMem_io_out_aluOp; // @[Core.scala 19:24]
  wire [2:0] ExRegMem_io_out_branch; // @[Core.scala 19:24]
  wire [1:0] ExRegMem_io_out_memtoReg; // @[Core.scala 19:24]
  wire  ExRegMem_io_out_memWr; // @[Core.scala 19:24]
  wire [2:0] ExRegMem_io_out_memOp; // @[Core.scala 19:24]
  wire  ExRegMem_io_out_rdEn; // @[Core.scala 19:24]
  wire [4:0] ExRegMem_io_out_rdAddr; // @[Core.scala 19:24]
  wire [63:0] ExRegMem_io_out_rs1Data; // @[Core.scala 19:24]
  wire [63:0] ExRegMem_io_out_rs2Data; // @[Core.scala 19:24]
  wire [63:0] ExRegMem_io_out_imm; // @[Core.scala 19:24]
  wire [63:0] ExRegMem_io_out_aluRes; // @[Core.scala 19:24]
  wire [63:0] ExRegMem_io_out_memData; // @[Core.scala 19:24]
  wire  ExRegMem_io_flush; // @[Core.scala 19:24]
  wire  ExRegMem_io_stall; // @[Core.scala 19:24]
  wire  MEM_clock; // @[Core.scala 20:19]
  wire  MEM_reset; // @[Core.scala 20:19]
  wire  MEM_io_dmem_data_valid; // @[Core.scala 20:19]
  wire  MEM_io_dmem_data_ready; // @[Core.scala 20:19]
  wire  MEM_io_dmem_data_req; // @[Core.scala 20:19]
  wire [31:0] MEM_io_dmem_data_addr; // @[Core.scala 20:19]
  wire [1:0] MEM_io_dmem_data_size; // @[Core.scala 20:19]
  wire [7:0] MEM_io_dmem_data_strb; // @[Core.scala 20:19]
  wire [63:0] MEM_io_dmem_data_read; // @[Core.scala 20:19]
  wire [127:0] MEM_io_dmem_data_write; // @[Core.scala 20:19]
  wire  MEM_io_in_valid; // @[Core.scala 20:19]
  wire [31:0] MEM_io_in_pc; // @[Core.scala 20:19]
  wire [31:0] MEM_io_in_inst; // @[Core.scala 20:19]
  wire  MEM_io_in_typeL; // @[Core.scala 20:19]
  wire  MEM_io_in_aluA; // @[Core.scala 20:19]
  wire [1:0] MEM_io_in_aluB; // @[Core.scala 20:19]
  wire [3:0] MEM_io_in_aluOp; // @[Core.scala 20:19]
  wire [2:0] MEM_io_in_branch; // @[Core.scala 20:19]
  wire [1:0] MEM_io_in_memtoReg; // @[Core.scala 20:19]
  wire  MEM_io_in_memWr; // @[Core.scala 20:19]
  wire [2:0] MEM_io_in_memOp; // @[Core.scala 20:19]
  wire  MEM_io_in_rdEn; // @[Core.scala 20:19]
  wire [4:0] MEM_io_in_rdAddr; // @[Core.scala 20:19]
  wire [63:0] MEM_io_in_rs1Data; // @[Core.scala 20:19]
  wire [63:0] MEM_io_in_rs2Data; // @[Core.scala 20:19]
  wire [63:0] MEM_io_in_imm; // @[Core.scala 20:19]
  wire [63:0] MEM_io_in_aluRes; // @[Core.scala 20:19]
  wire  MEM_io_out_valid; // @[Core.scala 20:19]
  wire [31:0] MEM_io_out_pc; // @[Core.scala 20:19]
  wire [31:0] MEM_io_out_inst; // @[Core.scala 20:19]
  wire  MEM_io_out_typeL; // @[Core.scala 20:19]
  wire  MEM_io_out_aluA; // @[Core.scala 20:19]
  wire [1:0] MEM_io_out_aluB; // @[Core.scala 20:19]
  wire [3:0] MEM_io_out_aluOp; // @[Core.scala 20:19]
  wire [2:0] MEM_io_out_branch; // @[Core.scala 20:19]
  wire [1:0] MEM_io_out_memtoReg; // @[Core.scala 20:19]
  wire  MEM_io_out_memWr; // @[Core.scala 20:19]
  wire [2:0] MEM_io_out_memOp; // @[Core.scala 20:19]
  wire  MEM_io_out_rdEn; // @[Core.scala 20:19]
  wire [4:0] MEM_io_out_rdAddr; // @[Core.scala 20:19]
  wire [63:0] MEM_io_out_rs1Data; // @[Core.scala 20:19]
  wire [63:0] MEM_io_out_rs2Data; // @[Core.scala 20:19]
  wire [63:0] MEM_io_out_imm; // @[Core.scala 20:19]
  wire [63:0] MEM_io_out_aluRes; // @[Core.scala 20:19]
  wire [63:0] MEM_io_out_memData; // @[Core.scala 20:19]
  wire  MEM_io_IFReady; // @[Core.scala 20:19]
  wire  MEM_io_memRdEn; // @[Core.scala 20:19]
  wire [4:0] MEM_io_memRdAddr; // @[Core.scala 20:19]
  wire [63:0] MEM_io_memRdData; // @[Core.scala 20:19]
  wire  MEM_io_memDone; // @[Core.scala 20:19]
  wire  MemRegWb_clock; // @[Core.scala 21:24]
  wire  MemRegWb_reset; // @[Core.scala 21:24]
  wire  MemRegWb_io_in_valid; // @[Core.scala 21:24]
  wire [31:0] MemRegWb_io_in_pc; // @[Core.scala 21:24]
  wire [31:0] MemRegWb_io_in_inst; // @[Core.scala 21:24]
  wire  MemRegWb_io_in_typeL; // @[Core.scala 21:24]
  wire  MemRegWb_io_in_aluA; // @[Core.scala 21:24]
  wire [1:0] MemRegWb_io_in_aluB; // @[Core.scala 21:24]
  wire [3:0] MemRegWb_io_in_aluOp; // @[Core.scala 21:24]
  wire [2:0] MemRegWb_io_in_branch; // @[Core.scala 21:24]
  wire [1:0] MemRegWb_io_in_memtoReg; // @[Core.scala 21:24]
  wire  MemRegWb_io_in_memWr; // @[Core.scala 21:24]
  wire [2:0] MemRegWb_io_in_memOp; // @[Core.scala 21:24]
  wire  MemRegWb_io_in_rdEn; // @[Core.scala 21:24]
  wire [4:0] MemRegWb_io_in_rdAddr; // @[Core.scala 21:24]
  wire [63:0] MemRegWb_io_in_rs1Data; // @[Core.scala 21:24]
  wire [63:0] MemRegWb_io_in_rs2Data; // @[Core.scala 21:24]
  wire [63:0] MemRegWb_io_in_imm; // @[Core.scala 21:24]
  wire [63:0] MemRegWb_io_in_aluRes; // @[Core.scala 21:24]
  wire [63:0] MemRegWb_io_in_memData; // @[Core.scala 21:24]
  wire  MemRegWb_io_out_valid; // @[Core.scala 21:24]
  wire [31:0] MemRegWb_io_out_pc; // @[Core.scala 21:24]
  wire [31:0] MemRegWb_io_out_inst; // @[Core.scala 21:24]
  wire  MemRegWb_io_out_typeL; // @[Core.scala 21:24]
  wire  MemRegWb_io_out_aluA; // @[Core.scala 21:24]
  wire [1:0] MemRegWb_io_out_aluB; // @[Core.scala 21:24]
  wire [3:0] MemRegWb_io_out_aluOp; // @[Core.scala 21:24]
  wire [2:0] MemRegWb_io_out_branch; // @[Core.scala 21:24]
  wire [1:0] MemRegWb_io_out_memtoReg; // @[Core.scala 21:24]
  wire  MemRegWb_io_out_memWr; // @[Core.scala 21:24]
  wire [2:0] MemRegWb_io_out_memOp; // @[Core.scala 21:24]
  wire  MemRegWb_io_out_rdEn; // @[Core.scala 21:24]
  wire [4:0] MemRegWb_io_out_rdAddr; // @[Core.scala 21:24]
  wire [63:0] MemRegWb_io_out_rs1Data; // @[Core.scala 21:24]
  wire [63:0] MemRegWb_io_out_rs2Data; // @[Core.scala 21:24]
  wire [63:0] MemRegWb_io_out_imm; // @[Core.scala 21:24]
  wire [63:0] MemRegWb_io_out_aluRes; // @[Core.scala 21:24]
  wire [63:0] MemRegWb_io_out_memData; // @[Core.scala 21:24]
  wire  MemRegWb_io_flush; // @[Core.scala 21:24]
  wire  MemRegWb_io_stall; // @[Core.scala 21:24]
  wire  WB_io_in_valid; // @[Core.scala 22:18]
  wire [31:0] WB_io_in_pc; // @[Core.scala 22:18]
  wire [31:0] WB_io_in_inst; // @[Core.scala 22:18]
  wire [1:0] WB_io_in_memtoReg; // @[Core.scala 22:18]
  wire  WB_io_in_rdEn; // @[Core.scala 22:18]
  wire [4:0] WB_io_in_rdAddr; // @[Core.scala 22:18]
  wire [63:0] WB_io_in_aluRes; // @[Core.scala 22:18]
  wire [63:0] WB_io_in_memData; // @[Core.scala 22:18]
  wire [31:0] WB_io_pc; // @[Core.scala 22:18]
  wire [31:0] WB_io_inst; // @[Core.scala 22:18]
  wire  WB_io_rdEn; // @[Core.scala 22:18]
  wire [4:0] WB_io_rdAddr; // @[Core.scala 22:18]
  wire [63:0] WB_io_rdData; // @[Core.scala 22:18]
  wire  WB_io_wbRdEn; // @[Core.scala 22:18]
  wire [4:0] WB_io_wbRdAddr; // @[Core.scala 22:18]
  wire [63:0] WB_io_wbRdData; // @[Core.scala 22:18]
  wire  WB_io_ready_cmt; // @[Core.scala 22:18]
  wire  dt_ic_clock; // @[Core.scala 103:21]
  wire [7:0] dt_ic_coreid; // @[Core.scala 103:21]
  wire [7:0] dt_ic_index; // @[Core.scala 103:21]
  wire  dt_ic_valid; // @[Core.scala 103:21]
  wire [63:0] dt_ic_pc; // @[Core.scala 103:21]
  wire [31:0] dt_ic_instr; // @[Core.scala 103:21]
  wire  dt_ic_skip; // @[Core.scala 103:21]
  wire  dt_ic_isRVC; // @[Core.scala 103:21]
  wire  dt_ic_scFailed; // @[Core.scala 103:21]
  wire  dt_ic_wen; // @[Core.scala 103:21]
  wire [63:0] dt_ic_wdata; // @[Core.scala 103:21]
  wire [7:0] dt_ic_wdest; // @[Core.scala 103:21]
  wire  dt_ae_clock; // @[Core.scala 117:21]
  wire [7:0] dt_ae_coreid; // @[Core.scala 117:21]
  wire [31:0] dt_ae_intrNO; // @[Core.scala 117:21]
  wire [31:0] dt_ae_cause; // @[Core.scala 117:21]
  wire [63:0] dt_ae_exceptionPC; // @[Core.scala 117:21]
  wire [31:0] dt_ae_exceptionInst; // @[Core.scala 117:21]
  wire  dt_te_clock; // @[Core.scala 133:21]
  wire [7:0] dt_te_coreid; // @[Core.scala 133:21]
  wire  dt_te_valid; // @[Core.scala 133:21]
  wire [2:0] dt_te_code; // @[Core.scala 133:21]
  wire [63:0] dt_te_pc; // @[Core.scala 133:21]
  wire [63:0] dt_te_cycleCnt; // @[Core.scala 133:21]
  wire [63:0] dt_te_instrCnt; // @[Core.scala 133:21]
  wire  dt_cs_clock; // @[Core.scala 142:21]
  wire [7:0] dt_cs_coreid; // @[Core.scala 142:21]
  wire [1:0] dt_cs_priviledgeMode; // @[Core.scala 142:21]
  wire [63:0] dt_cs_mstatus; // @[Core.scala 142:21]
  wire [63:0] dt_cs_sstatus; // @[Core.scala 142:21]
  wire [63:0] dt_cs_mepc; // @[Core.scala 142:21]
  wire [63:0] dt_cs_sepc; // @[Core.scala 142:21]
  wire [63:0] dt_cs_mtval; // @[Core.scala 142:21]
  wire [63:0] dt_cs_stval; // @[Core.scala 142:21]
  wire [63:0] dt_cs_mtvec; // @[Core.scala 142:21]
  wire [63:0] dt_cs_stvec; // @[Core.scala 142:21]
  wire [63:0] dt_cs_mcause; // @[Core.scala 142:21]
  wire [63:0] dt_cs_scause; // @[Core.scala 142:21]
  wire [63:0] dt_cs_satp; // @[Core.scala 142:21]
  wire [63:0] dt_cs_mip; // @[Core.scala 142:21]
  wire [63:0] dt_cs_mie; // @[Core.scala 142:21]
  wire [63:0] dt_cs_mscratch; // @[Core.scala 142:21]
  wire [63:0] dt_cs_sscratch; // @[Core.scala 142:21]
  wire [63:0] dt_cs_mideleg; // @[Core.scala 142:21]
  wire [63:0] dt_cs_medeleg; // @[Core.scala 142:21]
  wire  EXLHitID = ID_io_bubbleId & EX_io_bubbleEx; // @[Core.scala 25:33]
  wire  _flushIdExEn_T_1 = EX_io_pcSrc != 2'h0 | EXLHitID; // @[Core.scala 30:47]
  wire  valid = WB_io_ready_cmt & IF_io_IFDone & MEM_io_memDone; // @[Core.scala 101:47]
  reg  dt_ic_io_valid_REG; // @[Core.scala 107:31]
  reg [31:0] dt_ic_io_pc_REG; // @[Core.scala 108:31]
  reg [31:0] dt_ic_io_instr_REG; // @[Core.scala 109:31]
  reg  dt_ic_io_wen_REG; // @[Core.scala 113:31]
  reg [63:0] dt_ic_io_wdata_REG; // @[Core.scala 114:31]
  reg [4:0] dt_ic_io_wdest_REG; // @[Core.scala 115:31]
  reg [63:0] cycle_cnt; // @[Core.scala 124:26]
  reg [63:0] instr_cnt; // @[Core.scala 125:26]
  wire [63:0] _cycle_cnt_T_1 = cycle_cnt + 64'h1; // @[Core.scala 127:26]
  wire [63:0] _GEN_0 = {{63'd0}, valid}; // @[Core.scala 128:26]
  wire [63:0] _instr_cnt_T_1 = instr_cnt + _GEN_0; // @[Core.scala 128:26]
  wire [63:0] rf_a0_0 = ID_rf_10;
  InstFetch IF ( // @[Core.scala 14:18]
    .clock(IF_clock),
    .reset(IF_reset),
    .io_imem_inst_valid(IF_io_imem_inst_valid),
    .io_imem_inst_ready(IF_io_imem_inst_ready),
    .io_imem_inst_addr(IF_io_imem_inst_addr),
    .io_imem_inst_read(IF_io_imem_inst_read),
    .io_pcSrc(IF_io_pcSrc),
    .io_nextPC(IF_io_nextPC),
    .io_stall(IF_io_stall),
    .io_memDone(IF_io_memDone),
    .io_out_valid(IF_io_out_valid),
    .io_out_pc(IF_io_out_pc),
    .io_out_inst(IF_io_out_inst),
    .io_IFDone(IF_io_IFDone)
  );
  PipelineReg IfRegId ( // @[Core.scala 15:23]
    .clock(IfRegId_clock),
    .reset(IfRegId_reset),
    .io_in_valid(IfRegId_io_in_valid),
    .io_in_pc(IfRegId_io_in_pc),
    .io_in_inst(IfRegId_io_in_inst),
    .io_in_typeL(IfRegId_io_in_typeL),
    .io_in_aluA(IfRegId_io_in_aluA),
    .io_in_aluB(IfRegId_io_in_aluB),
    .io_in_aluOp(IfRegId_io_in_aluOp),
    .io_in_branch(IfRegId_io_in_branch),
    .io_in_memtoReg(IfRegId_io_in_memtoReg),
    .io_in_memWr(IfRegId_io_in_memWr),
    .io_in_memOp(IfRegId_io_in_memOp),
    .io_in_rdEn(IfRegId_io_in_rdEn),
    .io_in_rdAddr(IfRegId_io_in_rdAddr),
    .io_in_rs1Data(IfRegId_io_in_rs1Data),
    .io_in_rs2Data(IfRegId_io_in_rs2Data),
    .io_in_imm(IfRegId_io_in_imm),
    .io_in_aluRes(IfRegId_io_in_aluRes),
    .io_in_memData(IfRegId_io_in_memData),
    .io_out_valid(IfRegId_io_out_valid),
    .io_out_pc(IfRegId_io_out_pc),
    .io_out_inst(IfRegId_io_out_inst),
    .io_out_typeL(IfRegId_io_out_typeL),
    .io_out_aluA(IfRegId_io_out_aluA),
    .io_out_aluB(IfRegId_io_out_aluB),
    .io_out_aluOp(IfRegId_io_out_aluOp),
    .io_out_branch(IfRegId_io_out_branch),
    .io_out_memtoReg(IfRegId_io_out_memtoReg),
    .io_out_memWr(IfRegId_io_out_memWr),
    .io_out_memOp(IfRegId_io_out_memOp),
    .io_out_rdEn(IfRegId_io_out_rdEn),
    .io_out_rdAddr(IfRegId_io_out_rdAddr),
    .io_out_rs1Data(IfRegId_io_out_rs1Data),
    .io_out_rs2Data(IfRegId_io_out_rs2Data),
    .io_out_imm(IfRegId_io_out_imm),
    .io_out_aluRes(IfRegId_io_out_aluRes),
    .io_out_memData(IfRegId_io_out_memData),
    .io_flush(IfRegId_io_flush),
    .io_stall(IfRegId_io_stall)
  );
  Decode ID ( // @[Core.scala 16:18]
    .clock(ID_clock),
    .reset(ID_reset),
    .io_rdEn(ID_io_rdEn),
    .io_rdAddr(ID_io_rdAddr),
    .io_rdData(ID_io_rdData),
    .io_in_valid(ID_io_in_valid),
    .io_in_pc(ID_io_in_pc),
    .io_in_inst(ID_io_in_inst),
    .io_exeRdEn(ID_io_exeRdEn),
    .io_exeRdAddr(ID_io_exeRdAddr),
    .io_exeRdData(ID_io_exeRdData),
    .io_memRdEn(ID_io_memRdEn),
    .io_memRdAddr(ID_io_memRdAddr),
    .io_memRdData(ID_io_memRdData),
    .io_wbRdEn(ID_io_wbRdEn),
    .io_wbRdAddr(ID_io_wbRdAddr),
    .io_wbRdData(ID_io_wbRdData),
    .io_bubbleId(ID_io_bubbleId),
    .io_out_valid(ID_io_out_valid),
    .io_out_pc(ID_io_out_pc),
    .io_out_inst(ID_io_out_inst),
    .io_out_typeL(ID_io_out_typeL),
    .io_out_aluA(ID_io_out_aluA),
    .io_out_aluB(ID_io_out_aluB),
    .io_out_aluOp(ID_io_out_aluOp),
    .io_out_branch(ID_io_out_branch),
    .io_out_memtoReg(ID_io_out_memtoReg),
    .io_out_memWr(ID_io_out_memWr),
    .io_out_memOp(ID_io_out_memOp),
    .io_out_rdEn(ID_io_out_rdEn),
    .io_out_rdAddr(ID_io_out_rdAddr),
    .io_out_rs1Data(ID_io_out_rs1Data),
    .io_out_rs2Data(ID_io_out_rs2Data),
    .io_out_imm(ID_io_out_imm),
    .rf_10(ID_rf_10)
  );
  PipelineReg IdRegEx ( // @[Core.scala 17:23]
    .clock(IdRegEx_clock),
    .reset(IdRegEx_reset),
    .io_in_valid(IdRegEx_io_in_valid),
    .io_in_pc(IdRegEx_io_in_pc),
    .io_in_inst(IdRegEx_io_in_inst),
    .io_in_typeL(IdRegEx_io_in_typeL),
    .io_in_aluA(IdRegEx_io_in_aluA),
    .io_in_aluB(IdRegEx_io_in_aluB),
    .io_in_aluOp(IdRegEx_io_in_aluOp),
    .io_in_branch(IdRegEx_io_in_branch),
    .io_in_memtoReg(IdRegEx_io_in_memtoReg),
    .io_in_memWr(IdRegEx_io_in_memWr),
    .io_in_memOp(IdRegEx_io_in_memOp),
    .io_in_rdEn(IdRegEx_io_in_rdEn),
    .io_in_rdAddr(IdRegEx_io_in_rdAddr),
    .io_in_rs1Data(IdRegEx_io_in_rs1Data),
    .io_in_rs2Data(IdRegEx_io_in_rs2Data),
    .io_in_imm(IdRegEx_io_in_imm),
    .io_in_aluRes(IdRegEx_io_in_aluRes),
    .io_in_memData(IdRegEx_io_in_memData),
    .io_out_valid(IdRegEx_io_out_valid),
    .io_out_pc(IdRegEx_io_out_pc),
    .io_out_inst(IdRegEx_io_out_inst),
    .io_out_typeL(IdRegEx_io_out_typeL),
    .io_out_aluA(IdRegEx_io_out_aluA),
    .io_out_aluB(IdRegEx_io_out_aluB),
    .io_out_aluOp(IdRegEx_io_out_aluOp),
    .io_out_branch(IdRegEx_io_out_branch),
    .io_out_memtoReg(IdRegEx_io_out_memtoReg),
    .io_out_memWr(IdRegEx_io_out_memWr),
    .io_out_memOp(IdRegEx_io_out_memOp),
    .io_out_rdEn(IdRegEx_io_out_rdEn),
    .io_out_rdAddr(IdRegEx_io_out_rdAddr),
    .io_out_rs1Data(IdRegEx_io_out_rs1Data),
    .io_out_rs2Data(IdRegEx_io_out_rs2Data),
    .io_out_imm(IdRegEx_io_out_imm),
    .io_out_aluRes(IdRegEx_io_out_aluRes),
    .io_out_memData(IdRegEx_io_out_memData),
    .io_flush(IdRegEx_io_flush),
    .io_stall(IdRegEx_io_stall)
  );
  Execution EX ( // @[Core.scala 18:18]
    .io_in_valid(EX_io_in_valid),
    .io_in_pc(EX_io_in_pc),
    .io_in_inst(EX_io_in_inst),
    .io_in_typeL(EX_io_in_typeL),
    .io_in_aluA(EX_io_in_aluA),
    .io_in_aluB(EX_io_in_aluB),
    .io_in_aluOp(EX_io_in_aluOp),
    .io_in_branch(EX_io_in_branch),
    .io_in_memtoReg(EX_io_in_memtoReg),
    .io_in_memWr(EX_io_in_memWr),
    .io_in_memOp(EX_io_in_memOp),
    .io_in_rdEn(EX_io_in_rdEn),
    .io_in_rdAddr(EX_io_in_rdAddr),
    .io_in_rs1Data(EX_io_in_rs1Data),
    .io_in_rs2Data(EX_io_in_rs2Data),
    .io_in_imm(EX_io_in_imm),
    .io_out_valid(EX_io_out_valid),
    .io_out_pc(EX_io_out_pc),
    .io_out_inst(EX_io_out_inst),
    .io_out_typeL(EX_io_out_typeL),
    .io_out_aluA(EX_io_out_aluA),
    .io_out_aluB(EX_io_out_aluB),
    .io_out_aluOp(EX_io_out_aluOp),
    .io_out_branch(EX_io_out_branch),
    .io_out_memtoReg(EX_io_out_memtoReg),
    .io_out_memWr(EX_io_out_memWr),
    .io_out_memOp(EX_io_out_memOp),
    .io_out_rdEn(EX_io_out_rdEn),
    .io_out_rdAddr(EX_io_out_rdAddr),
    .io_out_rs1Data(EX_io_out_rs1Data),
    .io_out_rs2Data(EX_io_out_rs2Data),
    .io_out_imm(EX_io_out_imm),
    .io_out_aluRes(EX_io_out_aluRes),
    .io_exeRdEn(EX_io_exeRdEn),
    .io_exeRdAddr(EX_io_exeRdAddr),
    .io_exeRdData(EX_io_exeRdData),
    .io_bubbleEx(EX_io_bubbleEx),
    .io_pcSrc(EX_io_pcSrc),
    .io_nextPC(EX_io_nextPC)
  );
  PipelineReg ExRegMem ( // @[Core.scala 19:24]
    .clock(ExRegMem_clock),
    .reset(ExRegMem_reset),
    .io_in_valid(ExRegMem_io_in_valid),
    .io_in_pc(ExRegMem_io_in_pc),
    .io_in_inst(ExRegMem_io_in_inst),
    .io_in_typeL(ExRegMem_io_in_typeL),
    .io_in_aluA(ExRegMem_io_in_aluA),
    .io_in_aluB(ExRegMem_io_in_aluB),
    .io_in_aluOp(ExRegMem_io_in_aluOp),
    .io_in_branch(ExRegMem_io_in_branch),
    .io_in_memtoReg(ExRegMem_io_in_memtoReg),
    .io_in_memWr(ExRegMem_io_in_memWr),
    .io_in_memOp(ExRegMem_io_in_memOp),
    .io_in_rdEn(ExRegMem_io_in_rdEn),
    .io_in_rdAddr(ExRegMem_io_in_rdAddr),
    .io_in_rs1Data(ExRegMem_io_in_rs1Data),
    .io_in_rs2Data(ExRegMem_io_in_rs2Data),
    .io_in_imm(ExRegMem_io_in_imm),
    .io_in_aluRes(ExRegMem_io_in_aluRes),
    .io_in_memData(ExRegMem_io_in_memData),
    .io_out_valid(ExRegMem_io_out_valid),
    .io_out_pc(ExRegMem_io_out_pc),
    .io_out_inst(ExRegMem_io_out_inst),
    .io_out_typeL(ExRegMem_io_out_typeL),
    .io_out_aluA(ExRegMem_io_out_aluA),
    .io_out_aluB(ExRegMem_io_out_aluB),
    .io_out_aluOp(ExRegMem_io_out_aluOp),
    .io_out_branch(ExRegMem_io_out_branch),
    .io_out_memtoReg(ExRegMem_io_out_memtoReg),
    .io_out_memWr(ExRegMem_io_out_memWr),
    .io_out_memOp(ExRegMem_io_out_memOp),
    .io_out_rdEn(ExRegMem_io_out_rdEn),
    .io_out_rdAddr(ExRegMem_io_out_rdAddr),
    .io_out_rs1Data(ExRegMem_io_out_rs1Data),
    .io_out_rs2Data(ExRegMem_io_out_rs2Data),
    .io_out_imm(ExRegMem_io_out_imm),
    .io_out_aluRes(ExRegMem_io_out_aluRes),
    .io_out_memData(ExRegMem_io_out_memData),
    .io_flush(ExRegMem_io_flush),
    .io_stall(ExRegMem_io_stall)
  );
  DataMem MEM ( // @[Core.scala 20:19]
    .clock(MEM_clock),
    .reset(MEM_reset),
    .io_dmem_data_valid(MEM_io_dmem_data_valid),
    .io_dmem_data_ready(MEM_io_dmem_data_ready),
    .io_dmem_data_req(MEM_io_dmem_data_req),
    .io_dmem_data_addr(MEM_io_dmem_data_addr),
    .io_dmem_data_size(MEM_io_dmem_data_size),
    .io_dmem_data_strb(MEM_io_dmem_data_strb),
    .io_dmem_data_read(MEM_io_dmem_data_read),
    .io_dmem_data_write(MEM_io_dmem_data_write),
    .io_in_valid(MEM_io_in_valid),
    .io_in_pc(MEM_io_in_pc),
    .io_in_inst(MEM_io_in_inst),
    .io_in_typeL(MEM_io_in_typeL),
    .io_in_aluA(MEM_io_in_aluA),
    .io_in_aluB(MEM_io_in_aluB),
    .io_in_aluOp(MEM_io_in_aluOp),
    .io_in_branch(MEM_io_in_branch),
    .io_in_memtoReg(MEM_io_in_memtoReg),
    .io_in_memWr(MEM_io_in_memWr),
    .io_in_memOp(MEM_io_in_memOp),
    .io_in_rdEn(MEM_io_in_rdEn),
    .io_in_rdAddr(MEM_io_in_rdAddr),
    .io_in_rs1Data(MEM_io_in_rs1Data),
    .io_in_rs2Data(MEM_io_in_rs2Data),
    .io_in_imm(MEM_io_in_imm),
    .io_in_aluRes(MEM_io_in_aluRes),
    .io_out_valid(MEM_io_out_valid),
    .io_out_pc(MEM_io_out_pc),
    .io_out_inst(MEM_io_out_inst),
    .io_out_typeL(MEM_io_out_typeL),
    .io_out_aluA(MEM_io_out_aluA),
    .io_out_aluB(MEM_io_out_aluB),
    .io_out_aluOp(MEM_io_out_aluOp),
    .io_out_branch(MEM_io_out_branch),
    .io_out_memtoReg(MEM_io_out_memtoReg),
    .io_out_memWr(MEM_io_out_memWr),
    .io_out_memOp(MEM_io_out_memOp),
    .io_out_rdEn(MEM_io_out_rdEn),
    .io_out_rdAddr(MEM_io_out_rdAddr),
    .io_out_rs1Data(MEM_io_out_rs1Data),
    .io_out_rs2Data(MEM_io_out_rs2Data),
    .io_out_imm(MEM_io_out_imm),
    .io_out_aluRes(MEM_io_out_aluRes),
    .io_out_memData(MEM_io_out_memData),
    .io_IFReady(MEM_io_IFReady),
    .io_memRdEn(MEM_io_memRdEn),
    .io_memRdAddr(MEM_io_memRdAddr),
    .io_memRdData(MEM_io_memRdData),
    .io_memDone(MEM_io_memDone)
  );
  PipelineReg MemRegWb ( // @[Core.scala 21:24]
    .clock(MemRegWb_clock),
    .reset(MemRegWb_reset),
    .io_in_valid(MemRegWb_io_in_valid),
    .io_in_pc(MemRegWb_io_in_pc),
    .io_in_inst(MemRegWb_io_in_inst),
    .io_in_typeL(MemRegWb_io_in_typeL),
    .io_in_aluA(MemRegWb_io_in_aluA),
    .io_in_aluB(MemRegWb_io_in_aluB),
    .io_in_aluOp(MemRegWb_io_in_aluOp),
    .io_in_branch(MemRegWb_io_in_branch),
    .io_in_memtoReg(MemRegWb_io_in_memtoReg),
    .io_in_memWr(MemRegWb_io_in_memWr),
    .io_in_memOp(MemRegWb_io_in_memOp),
    .io_in_rdEn(MemRegWb_io_in_rdEn),
    .io_in_rdAddr(MemRegWb_io_in_rdAddr),
    .io_in_rs1Data(MemRegWb_io_in_rs1Data),
    .io_in_rs2Data(MemRegWb_io_in_rs2Data),
    .io_in_imm(MemRegWb_io_in_imm),
    .io_in_aluRes(MemRegWb_io_in_aluRes),
    .io_in_memData(MemRegWb_io_in_memData),
    .io_out_valid(MemRegWb_io_out_valid),
    .io_out_pc(MemRegWb_io_out_pc),
    .io_out_inst(MemRegWb_io_out_inst),
    .io_out_typeL(MemRegWb_io_out_typeL),
    .io_out_aluA(MemRegWb_io_out_aluA),
    .io_out_aluB(MemRegWb_io_out_aluB),
    .io_out_aluOp(MemRegWb_io_out_aluOp),
    .io_out_branch(MemRegWb_io_out_branch),
    .io_out_memtoReg(MemRegWb_io_out_memtoReg),
    .io_out_memWr(MemRegWb_io_out_memWr),
    .io_out_memOp(MemRegWb_io_out_memOp),
    .io_out_rdEn(MemRegWb_io_out_rdEn),
    .io_out_rdAddr(MemRegWb_io_out_rdAddr),
    .io_out_rs1Data(MemRegWb_io_out_rs1Data),
    .io_out_rs2Data(MemRegWb_io_out_rs2Data),
    .io_out_imm(MemRegWb_io_out_imm),
    .io_out_aluRes(MemRegWb_io_out_aluRes),
    .io_out_memData(MemRegWb_io_out_memData),
    .io_flush(MemRegWb_io_flush),
    .io_stall(MemRegWb_io_stall)
  );
  WriteBack WB ( // @[Core.scala 22:18]
    .io_in_valid(WB_io_in_valid),
    .io_in_pc(WB_io_in_pc),
    .io_in_inst(WB_io_in_inst),
    .io_in_memtoReg(WB_io_in_memtoReg),
    .io_in_rdEn(WB_io_in_rdEn),
    .io_in_rdAddr(WB_io_in_rdAddr),
    .io_in_aluRes(WB_io_in_aluRes),
    .io_in_memData(WB_io_in_memData),
    .io_pc(WB_io_pc),
    .io_inst(WB_io_inst),
    .io_rdEn(WB_io_rdEn),
    .io_rdAddr(WB_io_rdAddr),
    .io_rdData(WB_io_rdData),
    .io_wbRdEn(WB_io_wbRdEn),
    .io_wbRdAddr(WB_io_wbRdAddr),
    .io_wbRdData(WB_io_wbRdData),
    .io_ready_cmt(WB_io_ready_cmt)
  );
  DifftestInstrCommit dt_ic ( // @[Core.scala 103:21]
    .clock(dt_ic_clock),
    .coreid(dt_ic_coreid),
    .index(dt_ic_index),
    .valid(dt_ic_valid),
    .pc(dt_ic_pc),
    .instr(dt_ic_instr),
    .skip(dt_ic_skip),
    .isRVC(dt_ic_isRVC),
    .scFailed(dt_ic_scFailed),
    .wen(dt_ic_wen),
    .wdata(dt_ic_wdata),
    .wdest(dt_ic_wdest)
  );
  DifftestArchEvent dt_ae ( // @[Core.scala 117:21]
    .clock(dt_ae_clock),
    .coreid(dt_ae_coreid),
    .intrNO(dt_ae_intrNO),
    .cause(dt_ae_cause),
    .exceptionPC(dt_ae_exceptionPC),
    .exceptionInst(dt_ae_exceptionInst)
  );
  DifftestTrapEvent dt_te ( // @[Core.scala 133:21]
    .clock(dt_te_clock),
    .coreid(dt_te_coreid),
    .valid(dt_te_valid),
    .code(dt_te_code),
    .pc(dt_te_pc),
    .cycleCnt(dt_te_cycleCnt),
    .instrCnt(dt_te_instrCnt)
  );
  DifftestCSRState dt_cs ( // @[Core.scala 142:21]
    .clock(dt_cs_clock),
    .coreid(dt_cs_coreid),
    .priviledgeMode(dt_cs_priviledgeMode),
    .mstatus(dt_cs_mstatus),
    .sstatus(dt_cs_sstatus),
    .mepc(dt_cs_mepc),
    .sepc(dt_cs_sepc),
    .mtval(dt_cs_mtval),
    .stval(dt_cs_stval),
    .mtvec(dt_cs_mtvec),
    .stvec(dt_cs_stvec),
    .mcause(dt_cs_mcause),
    .scause(dt_cs_scause),
    .satp(dt_cs_satp),
    .mip(dt_cs_mip),
    .mie(dt_cs_mie),
    .mscratch(dt_cs_mscratch),
    .sscratch(dt_cs_sscratch),
    .mideleg(dt_cs_mideleg),
    .medeleg(dt_cs_medeleg)
  );
  assign io_imem_inst_valid = IF_io_imem_inst_valid; // @[Core.scala 47:22]
  assign io_imem_inst_addr = IF_io_imem_inst_addr; // @[Core.scala 49:21]
  assign io_dmem_data_valid = MEM_io_dmem_data_valid; // @[Core.scala 90:15]
  assign io_dmem_data_req = MEM_io_dmem_data_req; // @[Core.scala 90:15]
  assign io_dmem_data_addr = MEM_io_dmem_data_addr; // @[Core.scala 90:15]
  assign io_dmem_data_size = MEM_io_dmem_data_size; // @[Core.scala 90:15]
  assign io_dmem_data_strb = MEM_io_dmem_data_strb; // @[Core.scala 90:15]
  assign io_dmem_data_write = MEM_io_dmem_data_write; // @[Core.scala 90:15]
  assign IF_clock = clock;
  assign IF_reset = reset;
  assign IF_io_imem_inst_ready = io_imem_inst_ready; // @[Core.scala 53:25]
  assign IF_io_imem_inst_read = io_imem_inst_read; // @[Core.scala 52:24]
  assign IF_io_pcSrc = EX_io_pcSrc; // @[Core.scala 55:15]
  assign IF_io_nextPC = EX_io_nextPC; // @[Core.scala 56:16]
  assign IF_io_stall = EXLHitID | ~MEM_io_memDone; // @[Core.scala 57:27]
  assign IF_io_memDone = MEM_io_memDone; // @[Core.scala 58:17]
  assign IfRegId_clock = clock;
  assign IfRegId_reset = reset;
  assign IfRegId_io_in_valid = IF_io_out_valid; // @[Core.scala 60:17]
  assign IfRegId_io_in_pc = IF_io_out_pc; // @[Core.scala 60:17]
  assign IfRegId_io_in_inst = IF_io_out_inst; // @[Core.scala 60:17]
  assign IfRegId_io_in_typeL = 1'h0; // @[Core.scala 60:17]
  assign IfRegId_io_in_aluA = 1'h0; // @[Core.scala 60:17]
  assign IfRegId_io_in_aluB = 2'h0; // @[Core.scala 60:17]
  assign IfRegId_io_in_aluOp = 4'h0; // @[Core.scala 60:17]
  assign IfRegId_io_in_branch = 3'h0; // @[Core.scala 60:17]
  assign IfRegId_io_in_memtoReg = 2'h0; // @[Core.scala 60:17]
  assign IfRegId_io_in_memWr = 1'h0; // @[Core.scala 60:17]
  assign IfRegId_io_in_memOp = 3'h0; // @[Core.scala 60:17]
  assign IfRegId_io_in_rdEn = 1'h0; // @[Core.scala 60:17]
  assign IfRegId_io_in_rdAddr = 5'h0; // @[Core.scala 60:17]
  assign IfRegId_io_in_rs1Data = 64'h0; // @[Core.scala 60:17]
  assign IfRegId_io_in_rs2Data = 64'h0; // @[Core.scala 60:17]
  assign IfRegId_io_in_imm = 64'h0; // @[Core.scala 60:17]
  assign IfRegId_io_in_aluRes = 64'h0; // @[Core.scala 60:17]
  assign IfRegId_io_in_memData = 64'h0; // @[Core.scala 60:17]
  assign IfRegId_io_flush = 1'h0; // @[Core.scala 62:20]
  assign IfRegId_io_stall = ~IF_io_IFDone | EXLHitID; // @[Core.scala 39:36]
  assign ID_clock = clock;
  assign ID_reset = reset;
  assign ID_io_rdEn = WB_io_rdEn; // @[Core.scala 65:14]
  assign ID_io_rdAddr = WB_io_rdAddr; // @[Core.scala 66:16]
  assign ID_io_rdData = WB_io_rdData; // @[Core.scala 67:16]
  assign ID_io_in_valid = IfRegId_io_out_valid; // @[Core.scala 64:12]
  assign ID_io_in_pc = IfRegId_io_out_pc; // @[Core.scala 64:12]
  assign ID_io_in_inst = IfRegId_io_out_inst; // @[Core.scala 64:12]
  assign ID_io_exeRdEn = EX_io_exeRdEn; // @[Core.scala 69:17]
  assign ID_io_exeRdAddr = EX_io_exeRdAddr; // @[Core.scala 70:19]
  assign ID_io_exeRdData = EX_io_exeRdData; // @[Core.scala 71:19]
  assign ID_io_memRdEn = MEM_io_memRdEn; // @[Core.scala 72:17]
  assign ID_io_memRdAddr = MEM_io_memRdAddr; // @[Core.scala 73:19]
  assign ID_io_memRdData = MEM_io_memRdData; // @[Core.scala 74:19]
  assign ID_io_wbRdEn = WB_io_wbRdEn; // @[Core.scala 75:16]
  assign ID_io_wbRdAddr = WB_io_wbRdAddr; // @[Core.scala 76:18]
  assign ID_io_wbRdData = WB_io_wbRdData; // @[Core.scala 77:18]
  assign IdRegEx_clock = clock;
  assign IdRegEx_reset = reset;
  assign IdRegEx_io_in_valid = ID_io_out_valid; // @[Core.scala 79:17]
  assign IdRegEx_io_in_pc = ID_io_out_pc; // @[Core.scala 79:17]
  assign IdRegEx_io_in_inst = ID_io_out_inst; // @[Core.scala 79:17]
  assign IdRegEx_io_in_typeL = ID_io_out_typeL; // @[Core.scala 79:17]
  assign IdRegEx_io_in_aluA = ID_io_out_aluA; // @[Core.scala 79:17]
  assign IdRegEx_io_in_aluB = ID_io_out_aluB; // @[Core.scala 79:17]
  assign IdRegEx_io_in_aluOp = ID_io_out_aluOp; // @[Core.scala 79:17]
  assign IdRegEx_io_in_branch = ID_io_out_branch; // @[Core.scala 79:17]
  assign IdRegEx_io_in_memtoReg = ID_io_out_memtoReg; // @[Core.scala 79:17]
  assign IdRegEx_io_in_memWr = ID_io_out_memWr; // @[Core.scala 79:17]
  assign IdRegEx_io_in_memOp = ID_io_out_memOp; // @[Core.scala 79:17]
  assign IdRegEx_io_in_rdEn = ID_io_out_rdEn; // @[Core.scala 79:17]
  assign IdRegEx_io_in_rdAddr = ID_io_out_rdAddr; // @[Core.scala 79:17]
  assign IdRegEx_io_in_rs1Data = ID_io_out_rs1Data; // @[Core.scala 79:17]
  assign IdRegEx_io_in_rs2Data = ID_io_out_rs2Data; // @[Core.scala 79:17]
  assign IdRegEx_io_in_imm = ID_io_out_imm; // @[Core.scala 79:17]
  assign IdRegEx_io_in_aluRes = 64'h0; // @[Core.scala 79:17]
  assign IdRegEx_io_in_memData = 64'h0; // @[Core.scala 79:17]
  assign IdRegEx_io_flush = IF_io_IFDone & _flushIdExEn_T_1; // @[Core.scala 29:25]
  assign IdRegEx_io_stall = ~IF_io_IFDone; // @[Core.scala 40:22]
  assign EX_io_in_valid = IdRegEx_io_out_valid; // @[Core.scala 83:12]
  assign EX_io_in_pc = IdRegEx_io_out_pc; // @[Core.scala 83:12]
  assign EX_io_in_inst = IdRegEx_io_out_inst; // @[Core.scala 83:12]
  assign EX_io_in_typeL = IdRegEx_io_out_typeL; // @[Core.scala 83:12]
  assign EX_io_in_aluA = IdRegEx_io_out_aluA; // @[Core.scala 83:12]
  assign EX_io_in_aluB = IdRegEx_io_out_aluB; // @[Core.scala 83:12]
  assign EX_io_in_aluOp = IdRegEx_io_out_aluOp; // @[Core.scala 83:12]
  assign EX_io_in_branch = IdRegEx_io_out_branch; // @[Core.scala 83:12]
  assign EX_io_in_memtoReg = IdRegEx_io_out_memtoReg; // @[Core.scala 83:12]
  assign EX_io_in_memWr = IdRegEx_io_out_memWr; // @[Core.scala 83:12]
  assign EX_io_in_memOp = IdRegEx_io_out_memOp; // @[Core.scala 83:12]
  assign EX_io_in_rdEn = IdRegEx_io_out_rdEn; // @[Core.scala 83:12]
  assign EX_io_in_rdAddr = IdRegEx_io_out_rdAddr; // @[Core.scala 83:12]
  assign EX_io_in_rs1Data = IdRegEx_io_out_rs1Data; // @[Core.scala 83:12]
  assign EX_io_in_rs2Data = IdRegEx_io_out_rs2Data; // @[Core.scala 83:12]
  assign EX_io_in_imm = IdRegEx_io_out_imm; // @[Core.scala 83:12]
  assign ExRegMem_clock = clock;
  assign ExRegMem_reset = reset;
  assign ExRegMem_io_in_valid = EX_io_out_valid; // @[Core.scala 85:18]
  assign ExRegMem_io_in_pc = EX_io_out_pc; // @[Core.scala 85:18]
  assign ExRegMem_io_in_inst = EX_io_out_inst; // @[Core.scala 85:18]
  assign ExRegMem_io_in_typeL = EX_io_out_typeL; // @[Core.scala 85:18]
  assign ExRegMem_io_in_aluA = EX_io_out_aluA; // @[Core.scala 85:18]
  assign ExRegMem_io_in_aluB = EX_io_out_aluB; // @[Core.scala 85:18]
  assign ExRegMem_io_in_aluOp = EX_io_out_aluOp; // @[Core.scala 85:18]
  assign ExRegMem_io_in_branch = EX_io_out_branch; // @[Core.scala 85:18]
  assign ExRegMem_io_in_memtoReg = EX_io_out_memtoReg; // @[Core.scala 85:18]
  assign ExRegMem_io_in_memWr = EX_io_out_memWr; // @[Core.scala 85:18]
  assign ExRegMem_io_in_memOp = EX_io_out_memOp; // @[Core.scala 85:18]
  assign ExRegMem_io_in_rdEn = EX_io_out_rdEn; // @[Core.scala 85:18]
  assign ExRegMem_io_in_rdAddr = EX_io_out_rdAddr; // @[Core.scala 85:18]
  assign ExRegMem_io_in_rs1Data = EX_io_out_rs1Data; // @[Core.scala 85:18]
  assign ExRegMem_io_in_rs2Data = EX_io_out_rs2Data; // @[Core.scala 85:18]
  assign ExRegMem_io_in_imm = EX_io_out_imm; // @[Core.scala 85:18]
  assign ExRegMem_io_in_aluRes = EX_io_out_aluRes; // @[Core.scala 85:18]
  assign ExRegMem_io_in_memData = 64'h0; // @[Core.scala 85:18]
  assign ExRegMem_io_flush = 1'h0; // @[Core.scala 87:21]
  assign ExRegMem_io_stall = ~IF_io_IFDone; // @[Core.scala 41:22]
  assign MEM_clock = clock;
  assign MEM_reset = reset;
  assign MEM_io_dmem_data_ready = io_dmem_data_ready; // @[Core.scala 90:15]
  assign MEM_io_dmem_data_read = io_dmem_data_read; // @[Core.scala 90:15]
  assign MEM_io_in_valid = ExRegMem_io_out_valid; // @[Core.scala 89:13]
  assign MEM_io_in_pc = ExRegMem_io_out_pc; // @[Core.scala 89:13]
  assign MEM_io_in_inst = ExRegMem_io_out_inst; // @[Core.scala 89:13]
  assign MEM_io_in_typeL = ExRegMem_io_out_typeL; // @[Core.scala 89:13]
  assign MEM_io_in_aluA = ExRegMem_io_out_aluA; // @[Core.scala 89:13]
  assign MEM_io_in_aluB = ExRegMem_io_out_aluB; // @[Core.scala 89:13]
  assign MEM_io_in_aluOp = ExRegMem_io_out_aluOp; // @[Core.scala 89:13]
  assign MEM_io_in_branch = ExRegMem_io_out_branch; // @[Core.scala 89:13]
  assign MEM_io_in_memtoReg = ExRegMem_io_out_memtoReg; // @[Core.scala 89:13]
  assign MEM_io_in_memWr = ExRegMem_io_out_memWr; // @[Core.scala 89:13]
  assign MEM_io_in_memOp = ExRegMem_io_out_memOp; // @[Core.scala 89:13]
  assign MEM_io_in_rdEn = ExRegMem_io_out_rdEn; // @[Core.scala 89:13]
  assign MEM_io_in_rdAddr = ExRegMem_io_out_rdAddr; // @[Core.scala 89:13]
  assign MEM_io_in_rs1Data = ExRegMem_io_out_rs1Data; // @[Core.scala 89:13]
  assign MEM_io_in_rs2Data = ExRegMem_io_out_rs2Data; // @[Core.scala 89:13]
  assign MEM_io_in_imm = ExRegMem_io_out_imm; // @[Core.scala 89:13]
  assign MEM_io_in_aluRes = ExRegMem_io_out_aluRes; // @[Core.scala 89:13]
  assign MEM_io_IFReady = io_imem_inst_ready; // @[Core.scala 91:18]
  assign MemRegWb_clock = clock;
  assign MemRegWb_reset = reset;
  assign MemRegWb_io_in_valid = MEM_io_out_valid; // @[Core.scala 93:18]
  assign MemRegWb_io_in_pc = MEM_io_out_pc; // @[Core.scala 93:18]
  assign MemRegWb_io_in_inst = MEM_io_out_inst; // @[Core.scala 93:18]
  assign MemRegWb_io_in_typeL = MEM_io_out_typeL; // @[Core.scala 93:18]
  assign MemRegWb_io_in_aluA = MEM_io_out_aluA; // @[Core.scala 93:18]
  assign MemRegWb_io_in_aluB = MEM_io_out_aluB; // @[Core.scala 93:18]
  assign MemRegWb_io_in_aluOp = MEM_io_out_aluOp; // @[Core.scala 93:18]
  assign MemRegWb_io_in_branch = MEM_io_out_branch; // @[Core.scala 93:18]
  assign MemRegWb_io_in_memtoReg = MEM_io_out_memtoReg; // @[Core.scala 93:18]
  assign MemRegWb_io_in_memWr = MEM_io_out_memWr; // @[Core.scala 93:18]
  assign MemRegWb_io_in_memOp = MEM_io_out_memOp; // @[Core.scala 93:18]
  assign MemRegWb_io_in_rdEn = MEM_io_out_rdEn; // @[Core.scala 93:18]
  assign MemRegWb_io_in_rdAddr = MEM_io_out_rdAddr; // @[Core.scala 93:18]
  assign MemRegWb_io_in_rs1Data = MEM_io_out_rs1Data; // @[Core.scala 93:18]
  assign MemRegWb_io_in_rs2Data = MEM_io_out_rs2Data; // @[Core.scala 93:18]
  assign MemRegWb_io_in_imm = MEM_io_out_imm; // @[Core.scala 93:18]
  assign MemRegWb_io_in_aluRes = MEM_io_out_aluRes; // @[Core.scala 93:18]
  assign MemRegWb_io_in_memData = MEM_io_out_memData; // @[Core.scala 93:18]
  assign MemRegWb_io_flush = 1'h0; // @[Core.scala 95:21]
  assign MemRegWb_io_stall = ~IF_io_IFDone; // @[Core.scala 42:22]
  assign WB_io_in_valid = MemRegWb_io_out_valid; // @[Core.scala 97:12]
  assign WB_io_in_pc = MemRegWb_io_out_pc; // @[Core.scala 97:12]
  assign WB_io_in_inst = MemRegWb_io_out_inst; // @[Core.scala 97:12]
  assign WB_io_in_memtoReg = MemRegWb_io_out_memtoReg; // @[Core.scala 97:12]
  assign WB_io_in_rdEn = MemRegWb_io_out_rdEn; // @[Core.scala 97:12]
  assign WB_io_in_rdAddr = MemRegWb_io_out_rdAddr; // @[Core.scala 97:12]
  assign WB_io_in_aluRes = MemRegWb_io_out_aluRes; // @[Core.scala 97:12]
  assign WB_io_in_memData = MemRegWb_io_out_memData; // @[Core.scala 97:12]
  assign dt_ic_clock = clock; // @[Core.scala 104:21]
  assign dt_ic_coreid = 8'h0; // @[Core.scala 105:21]
  assign dt_ic_index = 8'h0; // @[Core.scala 106:21]
  assign dt_ic_valid = dt_ic_io_valid_REG; // @[Core.scala 107:21]
  assign dt_ic_pc = {{32'd0}, dt_ic_io_pc_REG}; // @[Core.scala 108:21]
  assign dt_ic_instr = dt_ic_io_instr_REG; // @[Core.scala 109:21]
  assign dt_ic_skip = 1'h0; // @[Core.scala 110:21]
  assign dt_ic_isRVC = 1'h0; // @[Core.scala 111:21]
  assign dt_ic_scFailed = 1'h0; // @[Core.scala 112:21]
  assign dt_ic_wen = dt_ic_io_wen_REG; // @[Core.scala 113:21]
  assign dt_ic_wdata = dt_ic_io_wdata_REG; // @[Core.scala 114:21]
  assign dt_ic_wdest = {{3'd0}, dt_ic_io_wdest_REG}; // @[Core.scala 115:21]
  assign dt_ae_clock = clock; // @[Core.scala 118:25]
  assign dt_ae_coreid = 8'h0; // @[Core.scala 119:25]
  assign dt_ae_intrNO = 32'h0; // @[Core.scala 120:25]
  assign dt_ae_cause = 32'h0; // @[Core.scala 121:25]
  assign dt_ae_exceptionPC = 64'h0; // @[Core.scala 122:25]
  assign dt_ae_exceptionInst = 32'h0;
  assign dt_te_clock = clock; // @[Core.scala 134:21]
  assign dt_te_coreid = 8'h0; // @[Core.scala 135:21]
  assign dt_te_valid = WB_io_inst == 32'h6b; // @[Core.scala 136:36]
  assign dt_te_code = rf_a0_0[2:0]; // @[Core.scala 137:29]
  assign dt_te_pc = {{32'd0}, WB_io_pc}; // @[Core.scala 138:21]
  assign dt_te_cycleCnt = cycle_cnt; // @[Core.scala 139:21]
  assign dt_te_instrCnt = instr_cnt; // @[Core.scala 140:21]
  assign dt_cs_clock = clock; // @[Core.scala 143:27]
  assign dt_cs_coreid = 8'h0; // @[Core.scala 144:27]
  assign dt_cs_priviledgeMode = 2'h3; // @[Core.scala 145:27]
  assign dt_cs_mstatus = 64'h0; // @[Core.scala 146:27]
  assign dt_cs_sstatus = 64'h0; // @[Core.scala 147:27]
  assign dt_cs_mepc = 64'h0; // @[Core.scala 148:27]
  assign dt_cs_sepc = 64'h0; // @[Core.scala 149:27]
  assign dt_cs_mtval = 64'h0; // @[Core.scala 150:27]
  assign dt_cs_stval = 64'h0; // @[Core.scala 151:27]
  assign dt_cs_mtvec = 64'h0; // @[Core.scala 152:27]
  assign dt_cs_stvec = 64'h0; // @[Core.scala 153:27]
  assign dt_cs_mcause = 64'h0; // @[Core.scala 154:27]
  assign dt_cs_scause = 64'h0; // @[Core.scala 155:27]
  assign dt_cs_satp = 64'h0; // @[Core.scala 156:27]
  assign dt_cs_mip = 64'h0; // @[Core.scala 157:27]
  assign dt_cs_mie = 64'h0; // @[Core.scala 158:27]
  assign dt_cs_mscratch = 64'h0; // @[Core.scala 159:27]
  assign dt_cs_sscratch = 64'h0; // @[Core.scala 160:27]
  assign dt_cs_mideleg = 64'h0; // @[Core.scala 161:27]
  assign dt_cs_medeleg = 64'h0; // @[Core.scala 162:27]
  always @(posedge clock) begin
    dt_ic_io_valid_REG <= WB_io_ready_cmt & IF_io_IFDone & MEM_io_memDone; // @[Core.scala 101:47]
    dt_ic_io_pc_REG <= WB_io_pc; // @[Core.scala 108:31]
    dt_ic_io_instr_REG <= WB_io_inst; // @[Core.scala 109:31]
    dt_ic_io_wen_REG <= WB_io_rdEn; // @[Core.scala 113:31]
    dt_ic_io_wdata_REG <= WB_io_rdData; // @[Core.scala 114:31]
    dt_ic_io_wdest_REG <= WB_io_rdAddr; // @[Core.scala 115:31]
    if (reset) begin // @[Core.scala 124:26]
      cycle_cnt <= 64'h0; // @[Core.scala 124:26]
    end else begin
      cycle_cnt <= _cycle_cnt_T_1; // @[Core.scala 127:13]
    end
    if (reset) begin // @[Core.scala 125:26]
      instr_cnt <= 64'h0; // @[Core.scala 125:26]
    end else begin
      instr_cnt <= _instr_cnt_T_1; // @[Core.scala 128:13]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  dt_ic_io_valid_REG = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  dt_ic_io_pc_REG = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  dt_ic_io_instr_REG = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  dt_ic_io_wen_REG = _RAND_3[0:0];
  _RAND_4 = {2{`RANDOM}};
  dt_ic_io_wdata_REG = _RAND_4[63:0];
  _RAND_5 = {1{`RANDOM}};
  dt_ic_io_wdest_REG = _RAND_5[4:0];
  _RAND_6 = {2{`RANDOM}};
  cycle_cnt = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  instr_cnt = _RAND_7[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ICache(
  input          clock,
  input          reset,
  input          io_imem_inst_valid,
  output         io_imem_inst_ready,
  input  [31:0]  io_imem_inst_addr,
  output [31:0]  io_imem_inst_read,
  output         io_out_inst_valid,
  input          io_out_inst_ready,
  output [31:0]  io_out_inst_addr,
  input  [127:0] io_out_inst_read
);
`ifdef RANDOMIZE_REG_INIT
  reg [127:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_645;
  reg [31:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_649;
  reg [31:0] _RAND_650;
  reg [31:0] _RAND_651;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
  reg [31:0] _RAND_654;
  reg [31:0] _RAND_655;
  reg [31:0] _RAND_656;
  reg [31:0] _RAND_657;
  reg [31:0] _RAND_658;
  reg [31:0] _RAND_659;
  reg [31:0] _RAND_660;
  reg [31:0] _RAND_661;
  reg [31:0] _RAND_662;
  reg [31:0] _RAND_663;
  reg [31:0] _RAND_664;
  reg [31:0] _RAND_665;
  reg [31:0] _RAND_666;
  reg [31:0] _RAND_667;
  reg [31:0] _RAND_668;
  reg [31:0] _RAND_669;
  reg [31:0] _RAND_670;
  reg [31:0] _RAND_671;
  reg [31:0] _RAND_672;
  reg [31:0] _RAND_673;
  reg [31:0] _RAND_674;
  reg [31:0] _RAND_675;
  reg [31:0] _RAND_676;
  reg [31:0] _RAND_677;
  reg [31:0] _RAND_678;
  reg [31:0] _RAND_679;
  reg [31:0] _RAND_680;
  reg [31:0] _RAND_681;
  reg [31:0] _RAND_682;
  reg [31:0] _RAND_683;
  reg [31:0] _RAND_684;
  reg [31:0] _RAND_685;
  reg [31:0] _RAND_686;
  reg [31:0] _RAND_687;
  reg [31:0] _RAND_688;
  reg [31:0] _RAND_689;
  reg [31:0] _RAND_690;
  reg [31:0] _RAND_691;
  reg [31:0] _RAND_692;
  reg [31:0] _RAND_693;
  reg [31:0] _RAND_694;
  reg [31:0] _RAND_695;
  reg [31:0] _RAND_696;
  reg [31:0] _RAND_697;
  reg [31:0] _RAND_698;
  reg [31:0] _RAND_699;
  reg [31:0] _RAND_700;
  reg [31:0] _RAND_701;
  reg [31:0] _RAND_702;
  reg [31:0] _RAND_703;
  reg [31:0] _RAND_704;
  reg [31:0] _RAND_705;
  reg [31:0] _RAND_706;
  reg [31:0] _RAND_707;
  reg [31:0] _RAND_708;
  reg [31:0] _RAND_709;
  reg [31:0] _RAND_710;
  reg [31:0] _RAND_711;
  reg [31:0] _RAND_712;
  reg [31:0] _RAND_713;
  reg [31:0] _RAND_714;
  reg [31:0] _RAND_715;
  reg [31:0] _RAND_716;
  reg [31:0] _RAND_717;
  reg [31:0] _RAND_718;
  reg [31:0] _RAND_719;
  reg [31:0] _RAND_720;
  reg [31:0] _RAND_721;
  reg [31:0] _RAND_722;
  reg [31:0] _RAND_723;
  reg [31:0] _RAND_724;
  reg [31:0] _RAND_725;
  reg [31:0] _RAND_726;
  reg [31:0] _RAND_727;
  reg [31:0] _RAND_728;
  reg [31:0] _RAND_729;
  reg [31:0] _RAND_730;
  reg [31:0] _RAND_731;
  reg [31:0] _RAND_732;
  reg [31:0] _RAND_733;
  reg [31:0] _RAND_734;
  reg [31:0] _RAND_735;
  reg [31:0] _RAND_736;
  reg [31:0] _RAND_737;
  reg [31:0] _RAND_738;
  reg [31:0] _RAND_739;
  reg [31:0] _RAND_740;
  reg [31:0] _RAND_741;
  reg [31:0] _RAND_742;
  reg [31:0] _RAND_743;
  reg [31:0] _RAND_744;
  reg [31:0] _RAND_745;
  reg [31:0] _RAND_746;
  reg [31:0] _RAND_747;
  reg [31:0] _RAND_748;
  reg [31:0] _RAND_749;
  reg [31:0] _RAND_750;
  reg [31:0] _RAND_751;
  reg [31:0] _RAND_752;
  reg [31:0] _RAND_753;
  reg [31:0] _RAND_754;
  reg [31:0] _RAND_755;
  reg [31:0] _RAND_756;
  reg [31:0] _RAND_757;
  reg [31:0] _RAND_758;
  reg [31:0] _RAND_759;
  reg [31:0] _RAND_760;
  reg [31:0] _RAND_761;
  reg [31:0] _RAND_762;
  reg [31:0] _RAND_763;
  reg [31:0] _RAND_764;
  reg [31:0] _RAND_765;
  reg [31:0] _RAND_766;
  reg [31:0] _RAND_767;
  reg [31:0] _RAND_768;
  reg [31:0] _RAND_769;
`endif // RANDOMIZE_REG_INIT
  wire [127:0] req_Q; // @[ICache.scala 51:19]
  wire  req_CLK; // @[ICache.scala 51:19]
  wire  req_CEN; // @[ICache.scala 51:19]
  wire  req_WEN; // @[ICache.scala 51:19]
  wire [7:0] req_A; // @[ICache.scala 51:19]
  wire [127:0] req_D; // @[ICache.scala 51:19]
  reg [127:0] cacheWData; // @[ICache.scala 22:27]
  reg  way0V_0; // @[ICache.scala 27:22]
  reg  way0V_1; // @[ICache.scala 27:22]
  reg  way0V_2; // @[ICache.scala 27:22]
  reg  way0V_3; // @[ICache.scala 27:22]
  reg  way0V_4; // @[ICache.scala 27:22]
  reg  way0V_5; // @[ICache.scala 27:22]
  reg  way0V_6; // @[ICache.scala 27:22]
  reg  way0V_7; // @[ICache.scala 27:22]
  reg  way0V_8; // @[ICache.scala 27:22]
  reg  way0V_9; // @[ICache.scala 27:22]
  reg  way0V_10; // @[ICache.scala 27:22]
  reg  way0V_11; // @[ICache.scala 27:22]
  reg  way0V_12; // @[ICache.scala 27:22]
  reg  way0V_13; // @[ICache.scala 27:22]
  reg  way0V_14; // @[ICache.scala 27:22]
  reg  way0V_15; // @[ICache.scala 27:22]
  reg  way0V_16; // @[ICache.scala 27:22]
  reg  way0V_17; // @[ICache.scala 27:22]
  reg  way0V_18; // @[ICache.scala 27:22]
  reg  way0V_19; // @[ICache.scala 27:22]
  reg  way0V_20; // @[ICache.scala 27:22]
  reg  way0V_21; // @[ICache.scala 27:22]
  reg  way0V_22; // @[ICache.scala 27:22]
  reg  way0V_23; // @[ICache.scala 27:22]
  reg  way0V_24; // @[ICache.scala 27:22]
  reg  way0V_25; // @[ICache.scala 27:22]
  reg  way0V_26; // @[ICache.scala 27:22]
  reg  way0V_27; // @[ICache.scala 27:22]
  reg  way0V_28; // @[ICache.scala 27:22]
  reg  way0V_29; // @[ICache.scala 27:22]
  reg  way0V_30; // @[ICache.scala 27:22]
  reg  way0V_31; // @[ICache.scala 27:22]
  reg  way0V_32; // @[ICache.scala 27:22]
  reg  way0V_33; // @[ICache.scala 27:22]
  reg  way0V_34; // @[ICache.scala 27:22]
  reg  way0V_35; // @[ICache.scala 27:22]
  reg  way0V_36; // @[ICache.scala 27:22]
  reg  way0V_37; // @[ICache.scala 27:22]
  reg  way0V_38; // @[ICache.scala 27:22]
  reg  way0V_39; // @[ICache.scala 27:22]
  reg  way0V_40; // @[ICache.scala 27:22]
  reg  way0V_41; // @[ICache.scala 27:22]
  reg  way0V_42; // @[ICache.scala 27:22]
  reg  way0V_43; // @[ICache.scala 27:22]
  reg  way0V_44; // @[ICache.scala 27:22]
  reg  way0V_45; // @[ICache.scala 27:22]
  reg  way0V_46; // @[ICache.scala 27:22]
  reg  way0V_47; // @[ICache.scala 27:22]
  reg  way0V_48; // @[ICache.scala 27:22]
  reg  way0V_49; // @[ICache.scala 27:22]
  reg  way0V_50; // @[ICache.scala 27:22]
  reg  way0V_51; // @[ICache.scala 27:22]
  reg  way0V_52; // @[ICache.scala 27:22]
  reg  way0V_53; // @[ICache.scala 27:22]
  reg  way0V_54; // @[ICache.scala 27:22]
  reg  way0V_55; // @[ICache.scala 27:22]
  reg  way0V_56; // @[ICache.scala 27:22]
  reg  way0V_57; // @[ICache.scala 27:22]
  reg  way0V_58; // @[ICache.scala 27:22]
  reg  way0V_59; // @[ICache.scala 27:22]
  reg  way0V_60; // @[ICache.scala 27:22]
  reg  way0V_61; // @[ICache.scala 27:22]
  reg  way0V_62; // @[ICache.scala 27:22]
  reg  way0V_63; // @[ICache.scala 27:22]
  reg  way0V_64; // @[ICache.scala 27:22]
  reg  way0V_65; // @[ICache.scala 27:22]
  reg  way0V_66; // @[ICache.scala 27:22]
  reg  way0V_67; // @[ICache.scala 27:22]
  reg  way0V_68; // @[ICache.scala 27:22]
  reg  way0V_69; // @[ICache.scala 27:22]
  reg  way0V_70; // @[ICache.scala 27:22]
  reg  way0V_71; // @[ICache.scala 27:22]
  reg  way0V_72; // @[ICache.scala 27:22]
  reg  way0V_73; // @[ICache.scala 27:22]
  reg  way0V_74; // @[ICache.scala 27:22]
  reg  way0V_75; // @[ICache.scala 27:22]
  reg  way0V_76; // @[ICache.scala 27:22]
  reg  way0V_77; // @[ICache.scala 27:22]
  reg  way0V_78; // @[ICache.scala 27:22]
  reg  way0V_79; // @[ICache.scala 27:22]
  reg  way0V_80; // @[ICache.scala 27:22]
  reg  way0V_81; // @[ICache.scala 27:22]
  reg  way0V_82; // @[ICache.scala 27:22]
  reg  way0V_83; // @[ICache.scala 27:22]
  reg  way0V_84; // @[ICache.scala 27:22]
  reg  way0V_85; // @[ICache.scala 27:22]
  reg  way0V_86; // @[ICache.scala 27:22]
  reg  way0V_87; // @[ICache.scala 27:22]
  reg  way0V_88; // @[ICache.scala 27:22]
  reg  way0V_89; // @[ICache.scala 27:22]
  reg  way0V_90; // @[ICache.scala 27:22]
  reg  way0V_91; // @[ICache.scala 27:22]
  reg  way0V_92; // @[ICache.scala 27:22]
  reg  way0V_93; // @[ICache.scala 27:22]
  reg  way0V_94; // @[ICache.scala 27:22]
  reg  way0V_95; // @[ICache.scala 27:22]
  reg  way0V_96; // @[ICache.scala 27:22]
  reg  way0V_97; // @[ICache.scala 27:22]
  reg  way0V_98; // @[ICache.scala 27:22]
  reg  way0V_99; // @[ICache.scala 27:22]
  reg  way0V_100; // @[ICache.scala 27:22]
  reg  way0V_101; // @[ICache.scala 27:22]
  reg  way0V_102; // @[ICache.scala 27:22]
  reg  way0V_103; // @[ICache.scala 27:22]
  reg  way0V_104; // @[ICache.scala 27:22]
  reg  way0V_105; // @[ICache.scala 27:22]
  reg  way0V_106; // @[ICache.scala 27:22]
  reg  way0V_107; // @[ICache.scala 27:22]
  reg  way0V_108; // @[ICache.scala 27:22]
  reg  way0V_109; // @[ICache.scala 27:22]
  reg  way0V_110; // @[ICache.scala 27:22]
  reg  way0V_111; // @[ICache.scala 27:22]
  reg  way0V_112; // @[ICache.scala 27:22]
  reg  way0V_113; // @[ICache.scala 27:22]
  reg  way0V_114; // @[ICache.scala 27:22]
  reg  way0V_115; // @[ICache.scala 27:22]
  reg  way0V_116; // @[ICache.scala 27:22]
  reg  way0V_117; // @[ICache.scala 27:22]
  reg  way0V_118; // @[ICache.scala 27:22]
  reg  way0V_119; // @[ICache.scala 27:22]
  reg  way0V_120; // @[ICache.scala 27:22]
  reg  way0V_121; // @[ICache.scala 27:22]
  reg  way0V_122; // @[ICache.scala 27:22]
  reg  way0V_123; // @[ICache.scala 27:22]
  reg  way0V_124; // @[ICache.scala 27:22]
  reg  way0V_125; // @[ICache.scala 27:22]
  reg  way0V_126; // @[ICache.scala 27:22]
  reg  way0V_127; // @[ICache.scala 27:22]
  reg [20:0] way0Tag_0; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_1; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_2; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_3; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_4; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_5; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_6; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_7; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_8; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_9; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_10; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_11; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_12; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_13; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_14; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_15; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_16; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_17; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_18; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_19; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_20; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_21; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_22; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_23; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_24; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_25; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_26; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_27; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_28; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_29; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_30; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_31; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_32; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_33; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_34; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_35; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_36; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_37; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_38; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_39; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_40; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_41; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_42; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_43; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_44; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_45; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_46; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_47; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_48; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_49; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_50; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_51; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_52; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_53; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_54; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_55; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_56; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_57; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_58; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_59; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_60; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_61; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_62; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_63; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_64; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_65; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_66; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_67; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_68; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_69; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_70; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_71; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_72; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_73; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_74; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_75; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_76; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_77; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_78; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_79; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_80; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_81; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_82; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_83; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_84; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_85; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_86; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_87; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_88; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_89; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_90; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_91; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_92; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_93; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_94; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_95; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_96; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_97; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_98; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_99; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_100; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_101; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_102; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_103; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_104; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_105; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_106; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_107; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_108; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_109; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_110; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_111; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_112; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_113; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_114; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_115; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_116; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_117; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_118; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_119; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_120; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_121; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_122; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_123; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_124; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_125; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_126; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_127; // @[ICache.scala 28:24]
  reg  way0Age_0; // @[ICache.scala 30:24]
  reg  way0Age_1; // @[ICache.scala 30:24]
  reg  way0Age_2; // @[ICache.scala 30:24]
  reg  way0Age_3; // @[ICache.scala 30:24]
  reg  way0Age_4; // @[ICache.scala 30:24]
  reg  way0Age_5; // @[ICache.scala 30:24]
  reg  way0Age_6; // @[ICache.scala 30:24]
  reg  way0Age_7; // @[ICache.scala 30:24]
  reg  way0Age_8; // @[ICache.scala 30:24]
  reg  way0Age_9; // @[ICache.scala 30:24]
  reg  way0Age_10; // @[ICache.scala 30:24]
  reg  way0Age_11; // @[ICache.scala 30:24]
  reg  way0Age_12; // @[ICache.scala 30:24]
  reg  way0Age_13; // @[ICache.scala 30:24]
  reg  way0Age_14; // @[ICache.scala 30:24]
  reg  way0Age_15; // @[ICache.scala 30:24]
  reg  way0Age_16; // @[ICache.scala 30:24]
  reg  way0Age_17; // @[ICache.scala 30:24]
  reg  way0Age_18; // @[ICache.scala 30:24]
  reg  way0Age_19; // @[ICache.scala 30:24]
  reg  way0Age_20; // @[ICache.scala 30:24]
  reg  way0Age_21; // @[ICache.scala 30:24]
  reg  way0Age_22; // @[ICache.scala 30:24]
  reg  way0Age_23; // @[ICache.scala 30:24]
  reg  way0Age_24; // @[ICache.scala 30:24]
  reg  way0Age_25; // @[ICache.scala 30:24]
  reg  way0Age_26; // @[ICache.scala 30:24]
  reg  way0Age_27; // @[ICache.scala 30:24]
  reg  way0Age_28; // @[ICache.scala 30:24]
  reg  way0Age_29; // @[ICache.scala 30:24]
  reg  way0Age_30; // @[ICache.scala 30:24]
  reg  way0Age_31; // @[ICache.scala 30:24]
  reg  way0Age_32; // @[ICache.scala 30:24]
  reg  way0Age_33; // @[ICache.scala 30:24]
  reg  way0Age_34; // @[ICache.scala 30:24]
  reg  way0Age_35; // @[ICache.scala 30:24]
  reg  way0Age_36; // @[ICache.scala 30:24]
  reg  way0Age_37; // @[ICache.scala 30:24]
  reg  way0Age_38; // @[ICache.scala 30:24]
  reg  way0Age_39; // @[ICache.scala 30:24]
  reg  way0Age_40; // @[ICache.scala 30:24]
  reg  way0Age_41; // @[ICache.scala 30:24]
  reg  way0Age_42; // @[ICache.scala 30:24]
  reg  way0Age_43; // @[ICache.scala 30:24]
  reg  way0Age_44; // @[ICache.scala 30:24]
  reg  way0Age_45; // @[ICache.scala 30:24]
  reg  way0Age_46; // @[ICache.scala 30:24]
  reg  way0Age_47; // @[ICache.scala 30:24]
  reg  way0Age_48; // @[ICache.scala 30:24]
  reg  way0Age_49; // @[ICache.scala 30:24]
  reg  way0Age_50; // @[ICache.scala 30:24]
  reg  way0Age_51; // @[ICache.scala 30:24]
  reg  way0Age_52; // @[ICache.scala 30:24]
  reg  way0Age_53; // @[ICache.scala 30:24]
  reg  way0Age_54; // @[ICache.scala 30:24]
  reg  way0Age_55; // @[ICache.scala 30:24]
  reg  way0Age_56; // @[ICache.scala 30:24]
  reg  way0Age_57; // @[ICache.scala 30:24]
  reg  way0Age_58; // @[ICache.scala 30:24]
  reg  way0Age_59; // @[ICache.scala 30:24]
  reg  way0Age_60; // @[ICache.scala 30:24]
  reg  way0Age_61; // @[ICache.scala 30:24]
  reg  way0Age_62; // @[ICache.scala 30:24]
  reg  way0Age_63; // @[ICache.scala 30:24]
  reg  way0Age_64; // @[ICache.scala 30:24]
  reg  way0Age_65; // @[ICache.scala 30:24]
  reg  way0Age_66; // @[ICache.scala 30:24]
  reg  way0Age_67; // @[ICache.scala 30:24]
  reg  way0Age_68; // @[ICache.scala 30:24]
  reg  way0Age_69; // @[ICache.scala 30:24]
  reg  way0Age_70; // @[ICache.scala 30:24]
  reg  way0Age_71; // @[ICache.scala 30:24]
  reg  way0Age_72; // @[ICache.scala 30:24]
  reg  way0Age_73; // @[ICache.scala 30:24]
  reg  way0Age_74; // @[ICache.scala 30:24]
  reg  way0Age_75; // @[ICache.scala 30:24]
  reg  way0Age_76; // @[ICache.scala 30:24]
  reg  way0Age_77; // @[ICache.scala 30:24]
  reg  way0Age_78; // @[ICache.scala 30:24]
  reg  way0Age_79; // @[ICache.scala 30:24]
  reg  way0Age_80; // @[ICache.scala 30:24]
  reg  way0Age_81; // @[ICache.scala 30:24]
  reg  way0Age_82; // @[ICache.scala 30:24]
  reg  way0Age_83; // @[ICache.scala 30:24]
  reg  way0Age_84; // @[ICache.scala 30:24]
  reg  way0Age_85; // @[ICache.scala 30:24]
  reg  way0Age_86; // @[ICache.scala 30:24]
  reg  way0Age_87; // @[ICache.scala 30:24]
  reg  way0Age_88; // @[ICache.scala 30:24]
  reg  way0Age_89; // @[ICache.scala 30:24]
  reg  way0Age_90; // @[ICache.scala 30:24]
  reg  way0Age_91; // @[ICache.scala 30:24]
  reg  way0Age_92; // @[ICache.scala 30:24]
  reg  way0Age_93; // @[ICache.scala 30:24]
  reg  way0Age_94; // @[ICache.scala 30:24]
  reg  way0Age_95; // @[ICache.scala 30:24]
  reg  way0Age_96; // @[ICache.scala 30:24]
  reg  way0Age_97; // @[ICache.scala 30:24]
  reg  way0Age_98; // @[ICache.scala 30:24]
  reg  way0Age_99; // @[ICache.scala 30:24]
  reg  way0Age_100; // @[ICache.scala 30:24]
  reg  way0Age_101; // @[ICache.scala 30:24]
  reg  way0Age_102; // @[ICache.scala 30:24]
  reg  way0Age_103; // @[ICache.scala 30:24]
  reg  way0Age_104; // @[ICache.scala 30:24]
  reg  way0Age_105; // @[ICache.scala 30:24]
  reg  way0Age_106; // @[ICache.scala 30:24]
  reg  way0Age_107; // @[ICache.scala 30:24]
  reg  way0Age_108; // @[ICache.scala 30:24]
  reg  way0Age_109; // @[ICache.scala 30:24]
  reg  way0Age_110; // @[ICache.scala 30:24]
  reg  way0Age_111; // @[ICache.scala 30:24]
  reg  way0Age_112; // @[ICache.scala 30:24]
  reg  way0Age_113; // @[ICache.scala 30:24]
  reg  way0Age_114; // @[ICache.scala 30:24]
  reg  way0Age_115; // @[ICache.scala 30:24]
  reg  way0Age_116; // @[ICache.scala 30:24]
  reg  way0Age_117; // @[ICache.scala 30:24]
  reg  way0Age_118; // @[ICache.scala 30:24]
  reg  way0Age_119; // @[ICache.scala 30:24]
  reg  way0Age_120; // @[ICache.scala 30:24]
  reg  way0Age_121; // @[ICache.scala 30:24]
  reg  way0Age_122; // @[ICache.scala 30:24]
  reg  way0Age_123; // @[ICache.scala 30:24]
  reg  way0Age_124; // @[ICache.scala 30:24]
  reg  way0Age_125; // @[ICache.scala 30:24]
  reg  way0Age_126; // @[ICache.scala 30:24]
  reg  way0Age_127; // @[ICache.scala 30:24]
  reg  way1V_0; // @[ICache.scala 32:22]
  reg  way1V_1; // @[ICache.scala 32:22]
  reg  way1V_2; // @[ICache.scala 32:22]
  reg  way1V_3; // @[ICache.scala 32:22]
  reg  way1V_4; // @[ICache.scala 32:22]
  reg  way1V_5; // @[ICache.scala 32:22]
  reg  way1V_6; // @[ICache.scala 32:22]
  reg  way1V_7; // @[ICache.scala 32:22]
  reg  way1V_8; // @[ICache.scala 32:22]
  reg  way1V_9; // @[ICache.scala 32:22]
  reg  way1V_10; // @[ICache.scala 32:22]
  reg  way1V_11; // @[ICache.scala 32:22]
  reg  way1V_12; // @[ICache.scala 32:22]
  reg  way1V_13; // @[ICache.scala 32:22]
  reg  way1V_14; // @[ICache.scala 32:22]
  reg  way1V_15; // @[ICache.scala 32:22]
  reg  way1V_16; // @[ICache.scala 32:22]
  reg  way1V_17; // @[ICache.scala 32:22]
  reg  way1V_18; // @[ICache.scala 32:22]
  reg  way1V_19; // @[ICache.scala 32:22]
  reg  way1V_20; // @[ICache.scala 32:22]
  reg  way1V_21; // @[ICache.scala 32:22]
  reg  way1V_22; // @[ICache.scala 32:22]
  reg  way1V_23; // @[ICache.scala 32:22]
  reg  way1V_24; // @[ICache.scala 32:22]
  reg  way1V_25; // @[ICache.scala 32:22]
  reg  way1V_26; // @[ICache.scala 32:22]
  reg  way1V_27; // @[ICache.scala 32:22]
  reg  way1V_28; // @[ICache.scala 32:22]
  reg  way1V_29; // @[ICache.scala 32:22]
  reg  way1V_30; // @[ICache.scala 32:22]
  reg  way1V_31; // @[ICache.scala 32:22]
  reg  way1V_32; // @[ICache.scala 32:22]
  reg  way1V_33; // @[ICache.scala 32:22]
  reg  way1V_34; // @[ICache.scala 32:22]
  reg  way1V_35; // @[ICache.scala 32:22]
  reg  way1V_36; // @[ICache.scala 32:22]
  reg  way1V_37; // @[ICache.scala 32:22]
  reg  way1V_38; // @[ICache.scala 32:22]
  reg  way1V_39; // @[ICache.scala 32:22]
  reg  way1V_40; // @[ICache.scala 32:22]
  reg  way1V_41; // @[ICache.scala 32:22]
  reg  way1V_42; // @[ICache.scala 32:22]
  reg  way1V_43; // @[ICache.scala 32:22]
  reg  way1V_44; // @[ICache.scala 32:22]
  reg  way1V_45; // @[ICache.scala 32:22]
  reg  way1V_46; // @[ICache.scala 32:22]
  reg  way1V_47; // @[ICache.scala 32:22]
  reg  way1V_48; // @[ICache.scala 32:22]
  reg  way1V_49; // @[ICache.scala 32:22]
  reg  way1V_50; // @[ICache.scala 32:22]
  reg  way1V_51; // @[ICache.scala 32:22]
  reg  way1V_52; // @[ICache.scala 32:22]
  reg  way1V_53; // @[ICache.scala 32:22]
  reg  way1V_54; // @[ICache.scala 32:22]
  reg  way1V_55; // @[ICache.scala 32:22]
  reg  way1V_56; // @[ICache.scala 32:22]
  reg  way1V_57; // @[ICache.scala 32:22]
  reg  way1V_58; // @[ICache.scala 32:22]
  reg  way1V_59; // @[ICache.scala 32:22]
  reg  way1V_60; // @[ICache.scala 32:22]
  reg  way1V_61; // @[ICache.scala 32:22]
  reg  way1V_62; // @[ICache.scala 32:22]
  reg  way1V_63; // @[ICache.scala 32:22]
  reg  way1V_64; // @[ICache.scala 32:22]
  reg  way1V_65; // @[ICache.scala 32:22]
  reg  way1V_66; // @[ICache.scala 32:22]
  reg  way1V_67; // @[ICache.scala 32:22]
  reg  way1V_68; // @[ICache.scala 32:22]
  reg  way1V_69; // @[ICache.scala 32:22]
  reg  way1V_70; // @[ICache.scala 32:22]
  reg  way1V_71; // @[ICache.scala 32:22]
  reg  way1V_72; // @[ICache.scala 32:22]
  reg  way1V_73; // @[ICache.scala 32:22]
  reg  way1V_74; // @[ICache.scala 32:22]
  reg  way1V_75; // @[ICache.scala 32:22]
  reg  way1V_76; // @[ICache.scala 32:22]
  reg  way1V_77; // @[ICache.scala 32:22]
  reg  way1V_78; // @[ICache.scala 32:22]
  reg  way1V_79; // @[ICache.scala 32:22]
  reg  way1V_80; // @[ICache.scala 32:22]
  reg  way1V_81; // @[ICache.scala 32:22]
  reg  way1V_82; // @[ICache.scala 32:22]
  reg  way1V_83; // @[ICache.scala 32:22]
  reg  way1V_84; // @[ICache.scala 32:22]
  reg  way1V_85; // @[ICache.scala 32:22]
  reg  way1V_86; // @[ICache.scala 32:22]
  reg  way1V_87; // @[ICache.scala 32:22]
  reg  way1V_88; // @[ICache.scala 32:22]
  reg  way1V_89; // @[ICache.scala 32:22]
  reg  way1V_90; // @[ICache.scala 32:22]
  reg  way1V_91; // @[ICache.scala 32:22]
  reg  way1V_92; // @[ICache.scala 32:22]
  reg  way1V_93; // @[ICache.scala 32:22]
  reg  way1V_94; // @[ICache.scala 32:22]
  reg  way1V_95; // @[ICache.scala 32:22]
  reg  way1V_96; // @[ICache.scala 32:22]
  reg  way1V_97; // @[ICache.scala 32:22]
  reg  way1V_98; // @[ICache.scala 32:22]
  reg  way1V_99; // @[ICache.scala 32:22]
  reg  way1V_100; // @[ICache.scala 32:22]
  reg  way1V_101; // @[ICache.scala 32:22]
  reg  way1V_102; // @[ICache.scala 32:22]
  reg  way1V_103; // @[ICache.scala 32:22]
  reg  way1V_104; // @[ICache.scala 32:22]
  reg  way1V_105; // @[ICache.scala 32:22]
  reg  way1V_106; // @[ICache.scala 32:22]
  reg  way1V_107; // @[ICache.scala 32:22]
  reg  way1V_108; // @[ICache.scala 32:22]
  reg  way1V_109; // @[ICache.scala 32:22]
  reg  way1V_110; // @[ICache.scala 32:22]
  reg  way1V_111; // @[ICache.scala 32:22]
  reg  way1V_112; // @[ICache.scala 32:22]
  reg  way1V_113; // @[ICache.scala 32:22]
  reg  way1V_114; // @[ICache.scala 32:22]
  reg  way1V_115; // @[ICache.scala 32:22]
  reg  way1V_116; // @[ICache.scala 32:22]
  reg  way1V_117; // @[ICache.scala 32:22]
  reg  way1V_118; // @[ICache.scala 32:22]
  reg  way1V_119; // @[ICache.scala 32:22]
  reg  way1V_120; // @[ICache.scala 32:22]
  reg  way1V_121; // @[ICache.scala 32:22]
  reg  way1V_122; // @[ICache.scala 32:22]
  reg  way1V_123; // @[ICache.scala 32:22]
  reg  way1V_124; // @[ICache.scala 32:22]
  reg  way1V_125; // @[ICache.scala 32:22]
  reg  way1V_126; // @[ICache.scala 32:22]
  reg  way1V_127; // @[ICache.scala 32:22]
  reg [20:0] way1Tag_0; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_1; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_2; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_3; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_4; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_5; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_6; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_7; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_8; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_9; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_10; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_11; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_12; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_13; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_14; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_15; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_16; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_17; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_18; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_19; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_20; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_21; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_22; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_23; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_24; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_25; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_26; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_27; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_28; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_29; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_30; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_31; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_32; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_33; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_34; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_35; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_36; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_37; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_38; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_39; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_40; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_41; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_42; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_43; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_44; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_45; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_46; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_47; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_48; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_49; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_50; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_51; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_52; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_53; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_54; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_55; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_56; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_57; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_58; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_59; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_60; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_61; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_62; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_63; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_64; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_65; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_66; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_67; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_68; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_69; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_70; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_71; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_72; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_73; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_74; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_75; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_76; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_77; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_78; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_79; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_80; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_81; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_82; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_83; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_84; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_85; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_86; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_87; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_88; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_89; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_90; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_91; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_92; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_93; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_94; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_95; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_96; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_97; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_98; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_99; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_100; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_101; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_102; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_103; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_104; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_105; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_106; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_107; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_108; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_109; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_110; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_111; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_112; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_113; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_114; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_115; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_116; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_117; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_118; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_119; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_120; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_121; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_122; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_123; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_124; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_125; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_126; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_127; // @[ICache.scala 33:24]
  reg  way1Age_0; // @[ICache.scala 35:24]
  reg  way1Age_1; // @[ICache.scala 35:24]
  reg  way1Age_2; // @[ICache.scala 35:24]
  reg  way1Age_3; // @[ICache.scala 35:24]
  reg  way1Age_4; // @[ICache.scala 35:24]
  reg  way1Age_5; // @[ICache.scala 35:24]
  reg  way1Age_6; // @[ICache.scala 35:24]
  reg  way1Age_7; // @[ICache.scala 35:24]
  reg  way1Age_8; // @[ICache.scala 35:24]
  reg  way1Age_9; // @[ICache.scala 35:24]
  reg  way1Age_10; // @[ICache.scala 35:24]
  reg  way1Age_11; // @[ICache.scala 35:24]
  reg  way1Age_12; // @[ICache.scala 35:24]
  reg  way1Age_13; // @[ICache.scala 35:24]
  reg  way1Age_14; // @[ICache.scala 35:24]
  reg  way1Age_15; // @[ICache.scala 35:24]
  reg  way1Age_16; // @[ICache.scala 35:24]
  reg  way1Age_17; // @[ICache.scala 35:24]
  reg  way1Age_18; // @[ICache.scala 35:24]
  reg  way1Age_19; // @[ICache.scala 35:24]
  reg  way1Age_20; // @[ICache.scala 35:24]
  reg  way1Age_21; // @[ICache.scala 35:24]
  reg  way1Age_22; // @[ICache.scala 35:24]
  reg  way1Age_23; // @[ICache.scala 35:24]
  reg  way1Age_24; // @[ICache.scala 35:24]
  reg  way1Age_25; // @[ICache.scala 35:24]
  reg  way1Age_26; // @[ICache.scala 35:24]
  reg  way1Age_27; // @[ICache.scala 35:24]
  reg  way1Age_28; // @[ICache.scala 35:24]
  reg  way1Age_29; // @[ICache.scala 35:24]
  reg  way1Age_30; // @[ICache.scala 35:24]
  reg  way1Age_31; // @[ICache.scala 35:24]
  reg  way1Age_32; // @[ICache.scala 35:24]
  reg  way1Age_33; // @[ICache.scala 35:24]
  reg  way1Age_34; // @[ICache.scala 35:24]
  reg  way1Age_35; // @[ICache.scala 35:24]
  reg  way1Age_36; // @[ICache.scala 35:24]
  reg  way1Age_37; // @[ICache.scala 35:24]
  reg  way1Age_38; // @[ICache.scala 35:24]
  reg  way1Age_39; // @[ICache.scala 35:24]
  reg  way1Age_40; // @[ICache.scala 35:24]
  reg  way1Age_41; // @[ICache.scala 35:24]
  reg  way1Age_42; // @[ICache.scala 35:24]
  reg  way1Age_43; // @[ICache.scala 35:24]
  reg  way1Age_44; // @[ICache.scala 35:24]
  reg  way1Age_45; // @[ICache.scala 35:24]
  reg  way1Age_46; // @[ICache.scala 35:24]
  reg  way1Age_47; // @[ICache.scala 35:24]
  reg  way1Age_48; // @[ICache.scala 35:24]
  reg  way1Age_49; // @[ICache.scala 35:24]
  reg  way1Age_50; // @[ICache.scala 35:24]
  reg  way1Age_51; // @[ICache.scala 35:24]
  reg  way1Age_52; // @[ICache.scala 35:24]
  reg  way1Age_53; // @[ICache.scala 35:24]
  reg  way1Age_54; // @[ICache.scala 35:24]
  reg  way1Age_55; // @[ICache.scala 35:24]
  reg  way1Age_56; // @[ICache.scala 35:24]
  reg  way1Age_57; // @[ICache.scala 35:24]
  reg  way1Age_58; // @[ICache.scala 35:24]
  reg  way1Age_59; // @[ICache.scala 35:24]
  reg  way1Age_60; // @[ICache.scala 35:24]
  reg  way1Age_61; // @[ICache.scala 35:24]
  reg  way1Age_62; // @[ICache.scala 35:24]
  reg  way1Age_63; // @[ICache.scala 35:24]
  reg  way1Age_64; // @[ICache.scala 35:24]
  reg  way1Age_65; // @[ICache.scala 35:24]
  reg  way1Age_66; // @[ICache.scala 35:24]
  reg  way1Age_67; // @[ICache.scala 35:24]
  reg  way1Age_68; // @[ICache.scala 35:24]
  reg  way1Age_69; // @[ICache.scala 35:24]
  reg  way1Age_70; // @[ICache.scala 35:24]
  reg  way1Age_71; // @[ICache.scala 35:24]
  reg  way1Age_72; // @[ICache.scala 35:24]
  reg  way1Age_73; // @[ICache.scala 35:24]
  reg  way1Age_74; // @[ICache.scala 35:24]
  reg  way1Age_75; // @[ICache.scala 35:24]
  reg  way1Age_76; // @[ICache.scala 35:24]
  reg  way1Age_77; // @[ICache.scala 35:24]
  reg  way1Age_78; // @[ICache.scala 35:24]
  reg  way1Age_79; // @[ICache.scala 35:24]
  reg  way1Age_80; // @[ICache.scala 35:24]
  reg  way1Age_81; // @[ICache.scala 35:24]
  reg  way1Age_82; // @[ICache.scala 35:24]
  reg  way1Age_83; // @[ICache.scala 35:24]
  reg  way1Age_84; // @[ICache.scala 35:24]
  reg  way1Age_85; // @[ICache.scala 35:24]
  reg  way1Age_86; // @[ICache.scala 35:24]
  reg  way1Age_87; // @[ICache.scala 35:24]
  reg  way1Age_88; // @[ICache.scala 35:24]
  reg  way1Age_89; // @[ICache.scala 35:24]
  reg  way1Age_90; // @[ICache.scala 35:24]
  reg  way1Age_91; // @[ICache.scala 35:24]
  reg  way1Age_92; // @[ICache.scala 35:24]
  reg  way1Age_93; // @[ICache.scala 35:24]
  reg  way1Age_94; // @[ICache.scala 35:24]
  reg  way1Age_95; // @[ICache.scala 35:24]
  reg  way1Age_96; // @[ICache.scala 35:24]
  reg  way1Age_97; // @[ICache.scala 35:24]
  reg  way1Age_98; // @[ICache.scala 35:24]
  reg  way1Age_99; // @[ICache.scala 35:24]
  reg  way1Age_100; // @[ICache.scala 35:24]
  reg  way1Age_101; // @[ICache.scala 35:24]
  reg  way1Age_102; // @[ICache.scala 35:24]
  reg  way1Age_103; // @[ICache.scala 35:24]
  reg  way1Age_104; // @[ICache.scala 35:24]
  reg  way1Age_105; // @[ICache.scala 35:24]
  reg  way1Age_106; // @[ICache.scala 35:24]
  reg  way1Age_107; // @[ICache.scala 35:24]
  reg  way1Age_108; // @[ICache.scala 35:24]
  reg  way1Age_109; // @[ICache.scala 35:24]
  reg  way1Age_110; // @[ICache.scala 35:24]
  reg  way1Age_111; // @[ICache.scala 35:24]
  reg  way1Age_112; // @[ICache.scala 35:24]
  reg  way1Age_113; // @[ICache.scala 35:24]
  reg  way1Age_114; // @[ICache.scala 35:24]
  reg  way1Age_115; // @[ICache.scala 35:24]
  reg  way1Age_116; // @[ICache.scala 35:24]
  reg  way1Age_117; // @[ICache.scala 35:24]
  reg  way1Age_118; // @[ICache.scala 35:24]
  reg  way1Age_119; // @[ICache.scala 35:24]
  reg  way1Age_120; // @[ICache.scala 35:24]
  reg  way1Age_121; // @[ICache.scala 35:24]
  reg  way1Age_122; // @[ICache.scala 35:24]
  reg  way1Age_123; // @[ICache.scala 35:24]
  reg  way1Age_124; // @[ICache.scala 35:24]
  reg  way1Age_125; // @[ICache.scala 35:24]
  reg  way1Age_126; // @[ICache.scala 35:24]
  reg  way1Age_127; // @[ICache.scala 35:24]
  reg [1:0] state; // @[ICache.scala 38:22]
  wire [20:0] reqTag = io_imem_inst_addr[31:11]; // @[ICache.scala 41:25]
  wire [6:0] reqIndex = io_imem_inst_addr[10:4]; // @[ICache.scala 42:27]
  wire [3:0] reqOff = io_imem_inst_addr[3:0]; // @[ICache.scala 43:25]
  wire [20:0] _GEN_1 = 7'h1 == reqIndex ? way0Tag_1 : way0Tag_0; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_2 = 7'h2 == reqIndex ? way0Tag_2 : _GEN_1; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_3 = 7'h3 == reqIndex ? way0Tag_3 : _GEN_2; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_4 = 7'h4 == reqIndex ? way0Tag_4 : _GEN_3; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_5 = 7'h5 == reqIndex ? way0Tag_5 : _GEN_4; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_6 = 7'h6 == reqIndex ? way0Tag_6 : _GEN_5; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_7 = 7'h7 == reqIndex ? way0Tag_7 : _GEN_6; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_8 = 7'h8 == reqIndex ? way0Tag_8 : _GEN_7; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_9 = 7'h9 == reqIndex ? way0Tag_9 : _GEN_8; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_10 = 7'ha == reqIndex ? way0Tag_10 : _GEN_9; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_11 = 7'hb == reqIndex ? way0Tag_11 : _GEN_10; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_12 = 7'hc == reqIndex ? way0Tag_12 : _GEN_11; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_13 = 7'hd == reqIndex ? way0Tag_13 : _GEN_12; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_14 = 7'he == reqIndex ? way0Tag_14 : _GEN_13; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_15 = 7'hf == reqIndex ? way0Tag_15 : _GEN_14; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_16 = 7'h10 == reqIndex ? way0Tag_16 : _GEN_15; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_17 = 7'h11 == reqIndex ? way0Tag_17 : _GEN_16; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_18 = 7'h12 == reqIndex ? way0Tag_18 : _GEN_17; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_19 = 7'h13 == reqIndex ? way0Tag_19 : _GEN_18; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_20 = 7'h14 == reqIndex ? way0Tag_20 : _GEN_19; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_21 = 7'h15 == reqIndex ? way0Tag_21 : _GEN_20; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_22 = 7'h16 == reqIndex ? way0Tag_22 : _GEN_21; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_23 = 7'h17 == reqIndex ? way0Tag_23 : _GEN_22; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_24 = 7'h18 == reqIndex ? way0Tag_24 : _GEN_23; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_25 = 7'h19 == reqIndex ? way0Tag_25 : _GEN_24; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_26 = 7'h1a == reqIndex ? way0Tag_26 : _GEN_25; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_27 = 7'h1b == reqIndex ? way0Tag_27 : _GEN_26; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_28 = 7'h1c == reqIndex ? way0Tag_28 : _GEN_27; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_29 = 7'h1d == reqIndex ? way0Tag_29 : _GEN_28; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_30 = 7'h1e == reqIndex ? way0Tag_30 : _GEN_29; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_31 = 7'h1f == reqIndex ? way0Tag_31 : _GEN_30; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_32 = 7'h20 == reqIndex ? way0Tag_32 : _GEN_31; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_33 = 7'h21 == reqIndex ? way0Tag_33 : _GEN_32; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_34 = 7'h22 == reqIndex ? way0Tag_34 : _GEN_33; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_35 = 7'h23 == reqIndex ? way0Tag_35 : _GEN_34; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_36 = 7'h24 == reqIndex ? way0Tag_36 : _GEN_35; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_37 = 7'h25 == reqIndex ? way0Tag_37 : _GEN_36; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_38 = 7'h26 == reqIndex ? way0Tag_38 : _GEN_37; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_39 = 7'h27 == reqIndex ? way0Tag_39 : _GEN_38; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_40 = 7'h28 == reqIndex ? way0Tag_40 : _GEN_39; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_41 = 7'h29 == reqIndex ? way0Tag_41 : _GEN_40; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_42 = 7'h2a == reqIndex ? way0Tag_42 : _GEN_41; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_43 = 7'h2b == reqIndex ? way0Tag_43 : _GEN_42; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_44 = 7'h2c == reqIndex ? way0Tag_44 : _GEN_43; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_45 = 7'h2d == reqIndex ? way0Tag_45 : _GEN_44; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_46 = 7'h2e == reqIndex ? way0Tag_46 : _GEN_45; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_47 = 7'h2f == reqIndex ? way0Tag_47 : _GEN_46; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_48 = 7'h30 == reqIndex ? way0Tag_48 : _GEN_47; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_49 = 7'h31 == reqIndex ? way0Tag_49 : _GEN_48; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_50 = 7'h32 == reqIndex ? way0Tag_50 : _GEN_49; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_51 = 7'h33 == reqIndex ? way0Tag_51 : _GEN_50; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_52 = 7'h34 == reqIndex ? way0Tag_52 : _GEN_51; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_53 = 7'h35 == reqIndex ? way0Tag_53 : _GEN_52; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_54 = 7'h36 == reqIndex ? way0Tag_54 : _GEN_53; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_55 = 7'h37 == reqIndex ? way0Tag_55 : _GEN_54; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_56 = 7'h38 == reqIndex ? way0Tag_56 : _GEN_55; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_57 = 7'h39 == reqIndex ? way0Tag_57 : _GEN_56; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_58 = 7'h3a == reqIndex ? way0Tag_58 : _GEN_57; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_59 = 7'h3b == reqIndex ? way0Tag_59 : _GEN_58; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_60 = 7'h3c == reqIndex ? way0Tag_60 : _GEN_59; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_61 = 7'h3d == reqIndex ? way0Tag_61 : _GEN_60; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_62 = 7'h3e == reqIndex ? way0Tag_62 : _GEN_61; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_63 = 7'h3f == reqIndex ? way0Tag_63 : _GEN_62; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_64 = 7'h40 == reqIndex ? way0Tag_64 : _GEN_63; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_65 = 7'h41 == reqIndex ? way0Tag_65 : _GEN_64; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_66 = 7'h42 == reqIndex ? way0Tag_66 : _GEN_65; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_67 = 7'h43 == reqIndex ? way0Tag_67 : _GEN_66; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_68 = 7'h44 == reqIndex ? way0Tag_68 : _GEN_67; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_69 = 7'h45 == reqIndex ? way0Tag_69 : _GEN_68; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_70 = 7'h46 == reqIndex ? way0Tag_70 : _GEN_69; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_71 = 7'h47 == reqIndex ? way0Tag_71 : _GEN_70; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_72 = 7'h48 == reqIndex ? way0Tag_72 : _GEN_71; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_73 = 7'h49 == reqIndex ? way0Tag_73 : _GEN_72; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_74 = 7'h4a == reqIndex ? way0Tag_74 : _GEN_73; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_75 = 7'h4b == reqIndex ? way0Tag_75 : _GEN_74; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_76 = 7'h4c == reqIndex ? way0Tag_76 : _GEN_75; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_77 = 7'h4d == reqIndex ? way0Tag_77 : _GEN_76; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_78 = 7'h4e == reqIndex ? way0Tag_78 : _GEN_77; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_79 = 7'h4f == reqIndex ? way0Tag_79 : _GEN_78; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_80 = 7'h50 == reqIndex ? way0Tag_80 : _GEN_79; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_81 = 7'h51 == reqIndex ? way0Tag_81 : _GEN_80; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_82 = 7'h52 == reqIndex ? way0Tag_82 : _GEN_81; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_83 = 7'h53 == reqIndex ? way0Tag_83 : _GEN_82; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_84 = 7'h54 == reqIndex ? way0Tag_84 : _GEN_83; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_85 = 7'h55 == reqIndex ? way0Tag_85 : _GEN_84; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_86 = 7'h56 == reqIndex ? way0Tag_86 : _GEN_85; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_87 = 7'h57 == reqIndex ? way0Tag_87 : _GEN_86; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_88 = 7'h58 == reqIndex ? way0Tag_88 : _GEN_87; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_89 = 7'h59 == reqIndex ? way0Tag_89 : _GEN_88; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_90 = 7'h5a == reqIndex ? way0Tag_90 : _GEN_89; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_91 = 7'h5b == reqIndex ? way0Tag_91 : _GEN_90; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_92 = 7'h5c == reqIndex ? way0Tag_92 : _GEN_91; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_93 = 7'h5d == reqIndex ? way0Tag_93 : _GEN_92; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_94 = 7'h5e == reqIndex ? way0Tag_94 : _GEN_93; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_95 = 7'h5f == reqIndex ? way0Tag_95 : _GEN_94; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_96 = 7'h60 == reqIndex ? way0Tag_96 : _GEN_95; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_97 = 7'h61 == reqIndex ? way0Tag_97 : _GEN_96; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_98 = 7'h62 == reqIndex ? way0Tag_98 : _GEN_97; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_99 = 7'h63 == reqIndex ? way0Tag_99 : _GEN_98; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_100 = 7'h64 == reqIndex ? way0Tag_100 : _GEN_99; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_101 = 7'h65 == reqIndex ? way0Tag_101 : _GEN_100; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_102 = 7'h66 == reqIndex ? way0Tag_102 : _GEN_101; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_103 = 7'h67 == reqIndex ? way0Tag_103 : _GEN_102; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_104 = 7'h68 == reqIndex ? way0Tag_104 : _GEN_103; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_105 = 7'h69 == reqIndex ? way0Tag_105 : _GEN_104; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_106 = 7'h6a == reqIndex ? way0Tag_106 : _GEN_105; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_107 = 7'h6b == reqIndex ? way0Tag_107 : _GEN_106; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_108 = 7'h6c == reqIndex ? way0Tag_108 : _GEN_107; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_109 = 7'h6d == reqIndex ? way0Tag_109 : _GEN_108; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_110 = 7'h6e == reqIndex ? way0Tag_110 : _GEN_109; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_111 = 7'h6f == reqIndex ? way0Tag_111 : _GEN_110; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_112 = 7'h70 == reqIndex ? way0Tag_112 : _GEN_111; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_113 = 7'h71 == reqIndex ? way0Tag_113 : _GEN_112; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_114 = 7'h72 == reqIndex ? way0Tag_114 : _GEN_113; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_115 = 7'h73 == reqIndex ? way0Tag_115 : _GEN_114; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_116 = 7'h74 == reqIndex ? way0Tag_116 : _GEN_115; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_117 = 7'h75 == reqIndex ? way0Tag_117 : _GEN_116; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_118 = 7'h76 == reqIndex ? way0Tag_118 : _GEN_117; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_119 = 7'h77 == reqIndex ? way0Tag_119 : _GEN_118; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_120 = 7'h78 == reqIndex ? way0Tag_120 : _GEN_119; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_121 = 7'h79 == reqIndex ? way0Tag_121 : _GEN_120; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_122 = 7'h7a == reqIndex ? way0Tag_122 : _GEN_121; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_123 = 7'h7b == reqIndex ? way0Tag_123 : _GEN_122; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_124 = 7'h7c == reqIndex ? way0Tag_124 : _GEN_123; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_125 = 7'h7d == reqIndex ? way0Tag_125 : _GEN_124; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_126 = 7'h7e == reqIndex ? way0Tag_126 : _GEN_125; // @[ICache.scala 45:{55,55}]
  wire [20:0] _GEN_127 = 7'h7f == reqIndex ? way0Tag_127 : _GEN_126; // @[ICache.scala 45:{55,55}]
  wire  _GEN_129 = 7'h1 == reqIndex ? way0V_1 : way0V_0; // @[ICache.scala 45:{33,33}]
  wire  _GEN_130 = 7'h2 == reqIndex ? way0V_2 : _GEN_129; // @[ICache.scala 45:{33,33}]
  wire  _GEN_131 = 7'h3 == reqIndex ? way0V_3 : _GEN_130; // @[ICache.scala 45:{33,33}]
  wire  _GEN_132 = 7'h4 == reqIndex ? way0V_4 : _GEN_131; // @[ICache.scala 45:{33,33}]
  wire  _GEN_133 = 7'h5 == reqIndex ? way0V_5 : _GEN_132; // @[ICache.scala 45:{33,33}]
  wire  _GEN_134 = 7'h6 == reqIndex ? way0V_6 : _GEN_133; // @[ICache.scala 45:{33,33}]
  wire  _GEN_135 = 7'h7 == reqIndex ? way0V_7 : _GEN_134; // @[ICache.scala 45:{33,33}]
  wire  _GEN_136 = 7'h8 == reqIndex ? way0V_8 : _GEN_135; // @[ICache.scala 45:{33,33}]
  wire  _GEN_137 = 7'h9 == reqIndex ? way0V_9 : _GEN_136; // @[ICache.scala 45:{33,33}]
  wire  _GEN_138 = 7'ha == reqIndex ? way0V_10 : _GEN_137; // @[ICache.scala 45:{33,33}]
  wire  _GEN_139 = 7'hb == reqIndex ? way0V_11 : _GEN_138; // @[ICache.scala 45:{33,33}]
  wire  _GEN_140 = 7'hc == reqIndex ? way0V_12 : _GEN_139; // @[ICache.scala 45:{33,33}]
  wire  _GEN_141 = 7'hd == reqIndex ? way0V_13 : _GEN_140; // @[ICache.scala 45:{33,33}]
  wire  _GEN_142 = 7'he == reqIndex ? way0V_14 : _GEN_141; // @[ICache.scala 45:{33,33}]
  wire  _GEN_143 = 7'hf == reqIndex ? way0V_15 : _GEN_142; // @[ICache.scala 45:{33,33}]
  wire  _GEN_144 = 7'h10 == reqIndex ? way0V_16 : _GEN_143; // @[ICache.scala 45:{33,33}]
  wire  _GEN_145 = 7'h11 == reqIndex ? way0V_17 : _GEN_144; // @[ICache.scala 45:{33,33}]
  wire  _GEN_146 = 7'h12 == reqIndex ? way0V_18 : _GEN_145; // @[ICache.scala 45:{33,33}]
  wire  _GEN_147 = 7'h13 == reqIndex ? way0V_19 : _GEN_146; // @[ICache.scala 45:{33,33}]
  wire  _GEN_148 = 7'h14 == reqIndex ? way0V_20 : _GEN_147; // @[ICache.scala 45:{33,33}]
  wire  _GEN_149 = 7'h15 == reqIndex ? way0V_21 : _GEN_148; // @[ICache.scala 45:{33,33}]
  wire  _GEN_150 = 7'h16 == reqIndex ? way0V_22 : _GEN_149; // @[ICache.scala 45:{33,33}]
  wire  _GEN_151 = 7'h17 == reqIndex ? way0V_23 : _GEN_150; // @[ICache.scala 45:{33,33}]
  wire  _GEN_152 = 7'h18 == reqIndex ? way0V_24 : _GEN_151; // @[ICache.scala 45:{33,33}]
  wire  _GEN_153 = 7'h19 == reqIndex ? way0V_25 : _GEN_152; // @[ICache.scala 45:{33,33}]
  wire  _GEN_154 = 7'h1a == reqIndex ? way0V_26 : _GEN_153; // @[ICache.scala 45:{33,33}]
  wire  _GEN_155 = 7'h1b == reqIndex ? way0V_27 : _GEN_154; // @[ICache.scala 45:{33,33}]
  wire  _GEN_156 = 7'h1c == reqIndex ? way0V_28 : _GEN_155; // @[ICache.scala 45:{33,33}]
  wire  _GEN_157 = 7'h1d == reqIndex ? way0V_29 : _GEN_156; // @[ICache.scala 45:{33,33}]
  wire  _GEN_158 = 7'h1e == reqIndex ? way0V_30 : _GEN_157; // @[ICache.scala 45:{33,33}]
  wire  _GEN_159 = 7'h1f == reqIndex ? way0V_31 : _GEN_158; // @[ICache.scala 45:{33,33}]
  wire  _GEN_160 = 7'h20 == reqIndex ? way0V_32 : _GEN_159; // @[ICache.scala 45:{33,33}]
  wire  _GEN_161 = 7'h21 == reqIndex ? way0V_33 : _GEN_160; // @[ICache.scala 45:{33,33}]
  wire  _GEN_162 = 7'h22 == reqIndex ? way0V_34 : _GEN_161; // @[ICache.scala 45:{33,33}]
  wire  _GEN_163 = 7'h23 == reqIndex ? way0V_35 : _GEN_162; // @[ICache.scala 45:{33,33}]
  wire  _GEN_164 = 7'h24 == reqIndex ? way0V_36 : _GEN_163; // @[ICache.scala 45:{33,33}]
  wire  _GEN_165 = 7'h25 == reqIndex ? way0V_37 : _GEN_164; // @[ICache.scala 45:{33,33}]
  wire  _GEN_166 = 7'h26 == reqIndex ? way0V_38 : _GEN_165; // @[ICache.scala 45:{33,33}]
  wire  _GEN_167 = 7'h27 == reqIndex ? way0V_39 : _GEN_166; // @[ICache.scala 45:{33,33}]
  wire  _GEN_168 = 7'h28 == reqIndex ? way0V_40 : _GEN_167; // @[ICache.scala 45:{33,33}]
  wire  _GEN_169 = 7'h29 == reqIndex ? way0V_41 : _GEN_168; // @[ICache.scala 45:{33,33}]
  wire  _GEN_170 = 7'h2a == reqIndex ? way0V_42 : _GEN_169; // @[ICache.scala 45:{33,33}]
  wire  _GEN_171 = 7'h2b == reqIndex ? way0V_43 : _GEN_170; // @[ICache.scala 45:{33,33}]
  wire  _GEN_172 = 7'h2c == reqIndex ? way0V_44 : _GEN_171; // @[ICache.scala 45:{33,33}]
  wire  _GEN_173 = 7'h2d == reqIndex ? way0V_45 : _GEN_172; // @[ICache.scala 45:{33,33}]
  wire  _GEN_174 = 7'h2e == reqIndex ? way0V_46 : _GEN_173; // @[ICache.scala 45:{33,33}]
  wire  _GEN_175 = 7'h2f == reqIndex ? way0V_47 : _GEN_174; // @[ICache.scala 45:{33,33}]
  wire  _GEN_176 = 7'h30 == reqIndex ? way0V_48 : _GEN_175; // @[ICache.scala 45:{33,33}]
  wire  _GEN_177 = 7'h31 == reqIndex ? way0V_49 : _GEN_176; // @[ICache.scala 45:{33,33}]
  wire  _GEN_178 = 7'h32 == reqIndex ? way0V_50 : _GEN_177; // @[ICache.scala 45:{33,33}]
  wire  _GEN_179 = 7'h33 == reqIndex ? way0V_51 : _GEN_178; // @[ICache.scala 45:{33,33}]
  wire  _GEN_180 = 7'h34 == reqIndex ? way0V_52 : _GEN_179; // @[ICache.scala 45:{33,33}]
  wire  _GEN_181 = 7'h35 == reqIndex ? way0V_53 : _GEN_180; // @[ICache.scala 45:{33,33}]
  wire  _GEN_182 = 7'h36 == reqIndex ? way0V_54 : _GEN_181; // @[ICache.scala 45:{33,33}]
  wire  _GEN_183 = 7'h37 == reqIndex ? way0V_55 : _GEN_182; // @[ICache.scala 45:{33,33}]
  wire  _GEN_184 = 7'h38 == reqIndex ? way0V_56 : _GEN_183; // @[ICache.scala 45:{33,33}]
  wire  _GEN_185 = 7'h39 == reqIndex ? way0V_57 : _GEN_184; // @[ICache.scala 45:{33,33}]
  wire  _GEN_186 = 7'h3a == reqIndex ? way0V_58 : _GEN_185; // @[ICache.scala 45:{33,33}]
  wire  _GEN_187 = 7'h3b == reqIndex ? way0V_59 : _GEN_186; // @[ICache.scala 45:{33,33}]
  wire  _GEN_188 = 7'h3c == reqIndex ? way0V_60 : _GEN_187; // @[ICache.scala 45:{33,33}]
  wire  _GEN_189 = 7'h3d == reqIndex ? way0V_61 : _GEN_188; // @[ICache.scala 45:{33,33}]
  wire  _GEN_190 = 7'h3e == reqIndex ? way0V_62 : _GEN_189; // @[ICache.scala 45:{33,33}]
  wire  _GEN_191 = 7'h3f == reqIndex ? way0V_63 : _GEN_190; // @[ICache.scala 45:{33,33}]
  wire  _GEN_192 = 7'h40 == reqIndex ? way0V_64 : _GEN_191; // @[ICache.scala 45:{33,33}]
  wire  _GEN_193 = 7'h41 == reqIndex ? way0V_65 : _GEN_192; // @[ICache.scala 45:{33,33}]
  wire  _GEN_194 = 7'h42 == reqIndex ? way0V_66 : _GEN_193; // @[ICache.scala 45:{33,33}]
  wire  _GEN_195 = 7'h43 == reqIndex ? way0V_67 : _GEN_194; // @[ICache.scala 45:{33,33}]
  wire  _GEN_196 = 7'h44 == reqIndex ? way0V_68 : _GEN_195; // @[ICache.scala 45:{33,33}]
  wire  _GEN_197 = 7'h45 == reqIndex ? way0V_69 : _GEN_196; // @[ICache.scala 45:{33,33}]
  wire  _GEN_198 = 7'h46 == reqIndex ? way0V_70 : _GEN_197; // @[ICache.scala 45:{33,33}]
  wire  _GEN_199 = 7'h47 == reqIndex ? way0V_71 : _GEN_198; // @[ICache.scala 45:{33,33}]
  wire  _GEN_200 = 7'h48 == reqIndex ? way0V_72 : _GEN_199; // @[ICache.scala 45:{33,33}]
  wire  _GEN_201 = 7'h49 == reqIndex ? way0V_73 : _GEN_200; // @[ICache.scala 45:{33,33}]
  wire  _GEN_202 = 7'h4a == reqIndex ? way0V_74 : _GEN_201; // @[ICache.scala 45:{33,33}]
  wire  _GEN_203 = 7'h4b == reqIndex ? way0V_75 : _GEN_202; // @[ICache.scala 45:{33,33}]
  wire  _GEN_204 = 7'h4c == reqIndex ? way0V_76 : _GEN_203; // @[ICache.scala 45:{33,33}]
  wire  _GEN_205 = 7'h4d == reqIndex ? way0V_77 : _GEN_204; // @[ICache.scala 45:{33,33}]
  wire  _GEN_206 = 7'h4e == reqIndex ? way0V_78 : _GEN_205; // @[ICache.scala 45:{33,33}]
  wire  _GEN_207 = 7'h4f == reqIndex ? way0V_79 : _GEN_206; // @[ICache.scala 45:{33,33}]
  wire  _GEN_208 = 7'h50 == reqIndex ? way0V_80 : _GEN_207; // @[ICache.scala 45:{33,33}]
  wire  _GEN_209 = 7'h51 == reqIndex ? way0V_81 : _GEN_208; // @[ICache.scala 45:{33,33}]
  wire  _GEN_210 = 7'h52 == reqIndex ? way0V_82 : _GEN_209; // @[ICache.scala 45:{33,33}]
  wire  _GEN_211 = 7'h53 == reqIndex ? way0V_83 : _GEN_210; // @[ICache.scala 45:{33,33}]
  wire  _GEN_212 = 7'h54 == reqIndex ? way0V_84 : _GEN_211; // @[ICache.scala 45:{33,33}]
  wire  _GEN_213 = 7'h55 == reqIndex ? way0V_85 : _GEN_212; // @[ICache.scala 45:{33,33}]
  wire  _GEN_214 = 7'h56 == reqIndex ? way0V_86 : _GEN_213; // @[ICache.scala 45:{33,33}]
  wire  _GEN_215 = 7'h57 == reqIndex ? way0V_87 : _GEN_214; // @[ICache.scala 45:{33,33}]
  wire  _GEN_216 = 7'h58 == reqIndex ? way0V_88 : _GEN_215; // @[ICache.scala 45:{33,33}]
  wire  _GEN_217 = 7'h59 == reqIndex ? way0V_89 : _GEN_216; // @[ICache.scala 45:{33,33}]
  wire  _GEN_218 = 7'h5a == reqIndex ? way0V_90 : _GEN_217; // @[ICache.scala 45:{33,33}]
  wire  _GEN_219 = 7'h5b == reqIndex ? way0V_91 : _GEN_218; // @[ICache.scala 45:{33,33}]
  wire  _GEN_220 = 7'h5c == reqIndex ? way0V_92 : _GEN_219; // @[ICache.scala 45:{33,33}]
  wire  _GEN_221 = 7'h5d == reqIndex ? way0V_93 : _GEN_220; // @[ICache.scala 45:{33,33}]
  wire  _GEN_222 = 7'h5e == reqIndex ? way0V_94 : _GEN_221; // @[ICache.scala 45:{33,33}]
  wire  _GEN_223 = 7'h5f == reqIndex ? way0V_95 : _GEN_222; // @[ICache.scala 45:{33,33}]
  wire  _GEN_224 = 7'h60 == reqIndex ? way0V_96 : _GEN_223; // @[ICache.scala 45:{33,33}]
  wire  _GEN_225 = 7'h61 == reqIndex ? way0V_97 : _GEN_224; // @[ICache.scala 45:{33,33}]
  wire  _GEN_226 = 7'h62 == reqIndex ? way0V_98 : _GEN_225; // @[ICache.scala 45:{33,33}]
  wire  _GEN_227 = 7'h63 == reqIndex ? way0V_99 : _GEN_226; // @[ICache.scala 45:{33,33}]
  wire  _GEN_228 = 7'h64 == reqIndex ? way0V_100 : _GEN_227; // @[ICache.scala 45:{33,33}]
  wire  _GEN_229 = 7'h65 == reqIndex ? way0V_101 : _GEN_228; // @[ICache.scala 45:{33,33}]
  wire  _GEN_230 = 7'h66 == reqIndex ? way0V_102 : _GEN_229; // @[ICache.scala 45:{33,33}]
  wire  _GEN_231 = 7'h67 == reqIndex ? way0V_103 : _GEN_230; // @[ICache.scala 45:{33,33}]
  wire  _GEN_232 = 7'h68 == reqIndex ? way0V_104 : _GEN_231; // @[ICache.scala 45:{33,33}]
  wire  _GEN_233 = 7'h69 == reqIndex ? way0V_105 : _GEN_232; // @[ICache.scala 45:{33,33}]
  wire  _GEN_234 = 7'h6a == reqIndex ? way0V_106 : _GEN_233; // @[ICache.scala 45:{33,33}]
  wire  _GEN_235 = 7'h6b == reqIndex ? way0V_107 : _GEN_234; // @[ICache.scala 45:{33,33}]
  wire  _GEN_236 = 7'h6c == reqIndex ? way0V_108 : _GEN_235; // @[ICache.scala 45:{33,33}]
  wire  _GEN_237 = 7'h6d == reqIndex ? way0V_109 : _GEN_236; // @[ICache.scala 45:{33,33}]
  wire  _GEN_238 = 7'h6e == reqIndex ? way0V_110 : _GEN_237; // @[ICache.scala 45:{33,33}]
  wire  _GEN_239 = 7'h6f == reqIndex ? way0V_111 : _GEN_238; // @[ICache.scala 45:{33,33}]
  wire  _GEN_240 = 7'h70 == reqIndex ? way0V_112 : _GEN_239; // @[ICache.scala 45:{33,33}]
  wire  _GEN_241 = 7'h71 == reqIndex ? way0V_113 : _GEN_240; // @[ICache.scala 45:{33,33}]
  wire  _GEN_242 = 7'h72 == reqIndex ? way0V_114 : _GEN_241; // @[ICache.scala 45:{33,33}]
  wire  _GEN_243 = 7'h73 == reqIndex ? way0V_115 : _GEN_242; // @[ICache.scala 45:{33,33}]
  wire  _GEN_244 = 7'h74 == reqIndex ? way0V_116 : _GEN_243; // @[ICache.scala 45:{33,33}]
  wire  _GEN_245 = 7'h75 == reqIndex ? way0V_117 : _GEN_244; // @[ICache.scala 45:{33,33}]
  wire  _GEN_246 = 7'h76 == reqIndex ? way0V_118 : _GEN_245; // @[ICache.scala 45:{33,33}]
  wire  _GEN_247 = 7'h77 == reqIndex ? way0V_119 : _GEN_246; // @[ICache.scala 45:{33,33}]
  wire  _GEN_248 = 7'h78 == reqIndex ? way0V_120 : _GEN_247; // @[ICache.scala 45:{33,33}]
  wire  _GEN_249 = 7'h79 == reqIndex ? way0V_121 : _GEN_248; // @[ICache.scala 45:{33,33}]
  wire  _GEN_250 = 7'h7a == reqIndex ? way0V_122 : _GEN_249; // @[ICache.scala 45:{33,33}]
  wire  _GEN_251 = 7'h7b == reqIndex ? way0V_123 : _GEN_250; // @[ICache.scala 45:{33,33}]
  wire  _GEN_252 = 7'h7c == reqIndex ? way0V_124 : _GEN_251; // @[ICache.scala 45:{33,33}]
  wire  _GEN_253 = 7'h7d == reqIndex ? way0V_125 : _GEN_252; // @[ICache.scala 45:{33,33}]
  wire  _GEN_254 = 7'h7e == reqIndex ? way0V_126 : _GEN_253; // @[ICache.scala 45:{33,33}]
  wire  _GEN_255 = 7'h7f == reqIndex ? way0V_127 : _GEN_254; // @[ICache.scala 45:{33,33}]
  wire  way0Hit = _GEN_255 & _GEN_127 == reqTag; // @[ICache.scala 45:33]
  wire [20:0] _GEN_257 = 7'h1 == reqIndex ? way1Tag_1 : way1Tag_0; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_258 = 7'h2 == reqIndex ? way1Tag_2 : _GEN_257; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_259 = 7'h3 == reqIndex ? way1Tag_3 : _GEN_258; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_260 = 7'h4 == reqIndex ? way1Tag_4 : _GEN_259; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_261 = 7'h5 == reqIndex ? way1Tag_5 : _GEN_260; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_262 = 7'h6 == reqIndex ? way1Tag_6 : _GEN_261; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_263 = 7'h7 == reqIndex ? way1Tag_7 : _GEN_262; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_264 = 7'h8 == reqIndex ? way1Tag_8 : _GEN_263; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_265 = 7'h9 == reqIndex ? way1Tag_9 : _GEN_264; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_266 = 7'ha == reqIndex ? way1Tag_10 : _GEN_265; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_267 = 7'hb == reqIndex ? way1Tag_11 : _GEN_266; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_268 = 7'hc == reqIndex ? way1Tag_12 : _GEN_267; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_269 = 7'hd == reqIndex ? way1Tag_13 : _GEN_268; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_270 = 7'he == reqIndex ? way1Tag_14 : _GEN_269; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_271 = 7'hf == reqIndex ? way1Tag_15 : _GEN_270; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_272 = 7'h10 == reqIndex ? way1Tag_16 : _GEN_271; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_273 = 7'h11 == reqIndex ? way1Tag_17 : _GEN_272; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_274 = 7'h12 == reqIndex ? way1Tag_18 : _GEN_273; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_275 = 7'h13 == reqIndex ? way1Tag_19 : _GEN_274; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_276 = 7'h14 == reqIndex ? way1Tag_20 : _GEN_275; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_277 = 7'h15 == reqIndex ? way1Tag_21 : _GEN_276; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_278 = 7'h16 == reqIndex ? way1Tag_22 : _GEN_277; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_279 = 7'h17 == reqIndex ? way1Tag_23 : _GEN_278; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_280 = 7'h18 == reqIndex ? way1Tag_24 : _GEN_279; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_281 = 7'h19 == reqIndex ? way1Tag_25 : _GEN_280; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_282 = 7'h1a == reqIndex ? way1Tag_26 : _GEN_281; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_283 = 7'h1b == reqIndex ? way1Tag_27 : _GEN_282; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_284 = 7'h1c == reqIndex ? way1Tag_28 : _GEN_283; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_285 = 7'h1d == reqIndex ? way1Tag_29 : _GEN_284; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_286 = 7'h1e == reqIndex ? way1Tag_30 : _GEN_285; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_287 = 7'h1f == reqIndex ? way1Tag_31 : _GEN_286; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_288 = 7'h20 == reqIndex ? way1Tag_32 : _GEN_287; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_289 = 7'h21 == reqIndex ? way1Tag_33 : _GEN_288; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_290 = 7'h22 == reqIndex ? way1Tag_34 : _GEN_289; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_291 = 7'h23 == reqIndex ? way1Tag_35 : _GEN_290; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_292 = 7'h24 == reqIndex ? way1Tag_36 : _GEN_291; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_293 = 7'h25 == reqIndex ? way1Tag_37 : _GEN_292; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_294 = 7'h26 == reqIndex ? way1Tag_38 : _GEN_293; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_295 = 7'h27 == reqIndex ? way1Tag_39 : _GEN_294; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_296 = 7'h28 == reqIndex ? way1Tag_40 : _GEN_295; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_297 = 7'h29 == reqIndex ? way1Tag_41 : _GEN_296; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_298 = 7'h2a == reqIndex ? way1Tag_42 : _GEN_297; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_299 = 7'h2b == reqIndex ? way1Tag_43 : _GEN_298; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_300 = 7'h2c == reqIndex ? way1Tag_44 : _GEN_299; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_301 = 7'h2d == reqIndex ? way1Tag_45 : _GEN_300; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_302 = 7'h2e == reqIndex ? way1Tag_46 : _GEN_301; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_303 = 7'h2f == reqIndex ? way1Tag_47 : _GEN_302; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_304 = 7'h30 == reqIndex ? way1Tag_48 : _GEN_303; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_305 = 7'h31 == reqIndex ? way1Tag_49 : _GEN_304; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_306 = 7'h32 == reqIndex ? way1Tag_50 : _GEN_305; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_307 = 7'h33 == reqIndex ? way1Tag_51 : _GEN_306; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_308 = 7'h34 == reqIndex ? way1Tag_52 : _GEN_307; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_309 = 7'h35 == reqIndex ? way1Tag_53 : _GEN_308; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_310 = 7'h36 == reqIndex ? way1Tag_54 : _GEN_309; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_311 = 7'h37 == reqIndex ? way1Tag_55 : _GEN_310; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_312 = 7'h38 == reqIndex ? way1Tag_56 : _GEN_311; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_313 = 7'h39 == reqIndex ? way1Tag_57 : _GEN_312; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_314 = 7'h3a == reqIndex ? way1Tag_58 : _GEN_313; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_315 = 7'h3b == reqIndex ? way1Tag_59 : _GEN_314; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_316 = 7'h3c == reqIndex ? way1Tag_60 : _GEN_315; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_317 = 7'h3d == reqIndex ? way1Tag_61 : _GEN_316; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_318 = 7'h3e == reqIndex ? way1Tag_62 : _GEN_317; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_319 = 7'h3f == reqIndex ? way1Tag_63 : _GEN_318; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_320 = 7'h40 == reqIndex ? way1Tag_64 : _GEN_319; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_321 = 7'h41 == reqIndex ? way1Tag_65 : _GEN_320; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_322 = 7'h42 == reqIndex ? way1Tag_66 : _GEN_321; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_323 = 7'h43 == reqIndex ? way1Tag_67 : _GEN_322; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_324 = 7'h44 == reqIndex ? way1Tag_68 : _GEN_323; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_325 = 7'h45 == reqIndex ? way1Tag_69 : _GEN_324; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_326 = 7'h46 == reqIndex ? way1Tag_70 : _GEN_325; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_327 = 7'h47 == reqIndex ? way1Tag_71 : _GEN_326; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_328 = 7'h48 == reqIndex ? way1Tag_72 : _GEN_327; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_329 = 7'h49 == reqIndex ? way1Tag_73 : _GEN_328; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_330 = 7'h4a == reqIndex ? way1Tag_74 : _GEN_329; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_331 = 7'h4b == reqIndex ? way1Tag_75 : _GEN_330; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_332 = 7'h4c == reqIndex ? way1Tag_76 : _GEN_331; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_333 = 7'h4d == reqIndex ? way1Tag_77 : _GEN_332; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_334 = 7'h4e == reqIndex ? way1Tag_78 : _GEN_333; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_335 = 7'h4f == reqIndex ? way1Tag_79 : _GEN_334; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_336 = 7'h50 == reqIndex ? way1Tag_80 : _GEN_335; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_337 = 7'h51 == reqIndex ? way1Tag_81 : _GEN_336; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_338 = 7'h52 == reqIndex ? way1Tag_82 : _GEN_337; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_339 = 7'h53 == reqIndex ? way1Tag_83 : _GEN_338; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_340 = 7'h54 == reqIndex ? way1Tag_84 : _GEN_339; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_341 = 7'h55 == reqIndex ? way1Tag_85 : _GEN_340; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_342 = 7'h56 == reqIndex ? way1Tag_86 : _GEN_341; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_343 = 7'h57 == reqIndex ? way1Tag_87 : _GEN_342; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_344 = 7'h58 == reqIndex ? way1Tag_88 : _GEN_343; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_345 = 7'h59 == reqIndex ? way1Tag_89 : _GEN_344; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_346 = 7'h5a == reqIndex ? way1Tag_90 : _GEN_345; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_347 = 7'h5b == reqIndex ? way1Tag_91 : _GEN_346; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_348 = 7'h5c == reqIndex ? way1Tag_92 : _GEN_347; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_349 = 7'h5d == reqIndex ? way1Tag_93 : _GEN_348; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_350 = 7'h5e == reqIndex ? way1Tag_94 : _GEN_349; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_351 = 7'h5f == reqIndex ? way1Tag_95 : _GEN_350; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_352 = 7'h60 == reqIndex ? way1Tag_96 : _GEN_351; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_353 = 7'h61 == reqIndex ? way1Tag_97 : _GEN_352; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_354 = 7'h62 == reqIndex ? way1Tag_98 : _GEN_353; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_355 = 7'h63 == reqIndex ? way1Tag_99 : _GEN_354; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_356 = 7'h64 == reqIndex ? way1Tag_100 : _GEN_355; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_357 = 7'h65 == reqIndex ? way1Tag_101 : _GEN_356; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_358 = 7'h66 == reqIndex ? way1Tag_102 : _GEN_357; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_359 = 7'h67 == reqIndex ? way1Tag_103 : _GEN_358; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_360 = 7'h68 == reqIndex ? way1Tag_104 : _GEN_359; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_361 = 7'h69 == reqIndex ? way1Tag_105 : _GEN_360; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_362 = 7'h6a == reqIndex ? way1Tag_106 : _GEN_361; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_363 = 7'h6b == reqIndex ? way1Tag_107 : _GEN_362; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_364 = 7'h6c == reqIndex ? way1Tag_108 : _GEN_363; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_365 = 7'h6d == reqIndex ? way1Tag_109 : _GEN_364; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_366 = 7'h6e == reqIndex ? way1Tag_110 : _GEN_365; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_367 = 7'h6f == reqIndex ? way1Tag_111 : _GEN_366; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_368 = 7'h70 == reqIndex ? way1Tag_112 : _GEN_367; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_369 = 7'h71 == reqIndex ? way1Tag_113 : _GEN_368; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_370 = 7'h72 == reqIndex ? way1Tag_114 : _GEN_369; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_371 = 7'h73 == reqIndex ? way1Tag_115 : _GEN_370; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_372 = 7'h74 == reqIndex ? way1Tag_116 : _GEN_371; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_373 = 7'h75 == reqIndex ? way1Tag_117 : _GEN_372; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_374 = 7'h76 == reqIndex ? way1Tag_118 : _GEN_373; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_375 = 7'h77 == reqIndex ? way1Tag_119 : _GEN_374; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_376 = 7'h78 == reqIndex ? way1Tag_120 : _GEN_375; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_377 = 7'h79 == reqIndex ? way1Tag_121 : _GEN_376; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_378 = 7'h7a == reqIndex ? way1Tag_122 : _GEN_377; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_379 = 7'h7b == reqIndex ? way1Tag_123 : _GEN_378; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_380 = 7'h7c == reqIndex ? way1Tag_124 : _GEN_379; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_381 = 7'h7d == reqIndex ? way1Tag_125 : _GEN_380; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_382 = 7'h7e == reqIndex ? way1Tag_126 : _GEN_381; // @[ICache.scala 46:{55,55}]
  wire [20:0] _GEN_383 = 7'h7f == reqIndex ? way1Tag_127 : _GEN_382; // @[ICache.scala 46:{55,55}]
  wire  _GEN_385 = 7'h1 == reqIndex ? way1V_1 : way1V_0; // @[ICache.scala 46:{33,33}]
  wire  _GEN_386 = 7'h2 == reqIndex ? way1V_2 : _GEN_385; // @[ICache.scala 46:{33,33}]
  wire  _GEN_387 = 7'h3 == reqIndex ? way1V_3 : _GEN_386; // @[ICache.scala 46:{33,33}]
  wire  _GEN_388 = 7'h4 == reqIndex ? way1V_4 : _GEN_387; // @[ICache.scala 46:{33,33}]
  wire  _GEN_389 = 7'h5 == reqIndex ? way1V_5 : _GEN_388; // @[ICache.scala 46:{33,33}]
  wire  _GEN_390 = 7'h6 == reqIndex ? way1V_6 : _GEN_389; // @[ICache.scala 46:{33,33}]
  wire  _GEN_391 = 7'h7 == reqIndex ? way1V_7 : _GEN_390; // @[ICache.scala 46:{33,33}]
  wire  _GEN_392 = 7'h8 == reqIndex ? way1V_8 : _GEN_391; // @[ICache.scala 46:{33,33}]
  wire  _GEN_393 = 7'h9 == reqIndex ? way1V_9 : _GEN_392; // @[ICache.scala 46:{33,33}]
  wire  _GEN_394 = 7'ha == reqIndex ? way1V_10 : _GEN_393; // @[ICache.scala 46:{33,33}]
  wire  _GEN_395 = 7'hb == reqIndex ? way1V_11 : _GEN_394; // @[ICache.scala 46:{33,33}]
  wire  _GEN_396 = 7'hc == reqIndex ? way1V_12 : _GEN_395; // @[ICache.scala 46:{33,33}]
  wire  _GEN_397 = 7'hd == reqIndex ? way1V_13 : _GEN_396; // @[ICache.scala 46:{33,33}]
  wire  _GEN_398 = 7'he == reqIndex ? way1V_14 : _GEN_397; // @[ICache.scala 46:{33,33}]
  wire  _GEN_399 = 7'hf == reqIndex ? way1V_15 : _GEN_398; // @[ICache.scala 46:{33,33}]
  wire  _GEN_400 = 7'h10 == reqIndex ? way1V_16 : _GEN_399; // @[ICache.scala 46:{33,33}]
  wire  _GEN_401 = 7'h11 == reqIndex ? way1V_17 : _GEN_400; // @[ICache.scala 46:{33,33}]
  wire  _GEN_402 = 7'h12 == reqIndex ? way1V_18 : _GEN_401; // @[ICache.scala 46:{33,33}]
  wire  _GEN_403 = 7'h13 == reqIndex ? way1V_19 : _GEN_402; // @[ICache.scala 46:{33,33}]
  wire  _GEN_404 = 7'h14 == reqIndex ? way1V_20 : _GEN_403; // @[ICache.scala 46:{33,33}]
  wire  _GEN_405 = 7'h15 == reqIndex ? way1V_21 : _GEN_404; // @[ICache.scala 46:{33,33}]
  wire  _GEN_406 = 7'h16 == reqIndex ? way1V_22 : _GEN_405; // @[ICache.scala 46:{33,33}]
  wire  _GEN_407 = 7'h17 == reqIndex ? way1V_23 : _GEN_406; // @[ICache.scala 46:{33,33}]
  wire  _GEN_408 = 7'h18 == reqIndex ? way1V_24 : _GEN_407; // @[ICache.scala 46:{33,33}]
  wire  _GEN_409 = 7'h19 == reqIndex ? way1V_25 : _GEN_408; // @[ICache.scala 46:{33,33}]
  wire  _GEN_410 = 7'h1a == reqIndex ? way1V_26 : _GEN_409; // @[ICache.scala 46:{33,33}]
  wire  _GEN_411 = 7'h1b == reqIndex ? way1V_27 : _GEN_410; // @[ICache.scala 46:{33,33}]
  wire  _GEN_412 = 7'h1c == reqIndex ? way1V_28 : _GEN_411; // @[ICache.scala 46:{33,33}]
  wire  _GEN_413 = 7'h1d == reqIndex ? way1V_29 : _GEN_412; // @[ICache.scala 46:{33,33}]
  wire  _GEN_414 = 7'h1e == reqIndex ? way1V_30 : _GEN_413; // @[ICache.scala 46:{33,33}]
  wire  _GEN_415 = 7'h1f == reqIndex ? way1V_31 : _GEN_414; // @[ICache.scala 46:{33,33}]
  wire  _GEN_416 = 7'h20 == reqIndex ? way1V_32 : _GEN_415; // @[ICache.scala 46:{33,33}]
  wire  _GEN_417 = 7'h21 == reqIndex ? way1V_33 : _GEN_416; // @[ICache.scala 46:{33,33}]
  wire  _GEN_418 = 7'h22 == reqIndex ? way1V_34 : _GEN_417; // @[ICache.scala 46:{33,33}]
  wire  _GEN_419 = 7'h23 == reqIndex ? way1V_35 : _GEN_418; // @[ICache.scala 46:{33,33}]
  wire  _GEN_420 = 7'h24 == reqIndex ? way1V_36 : _GEN_419; // @[ICache.scala 46:{33,33}]
  wire  _GEN_421 = 7'h25 == reqIndex ? way1V_37 : _GEN_420; // @[ICache.scala 46:{33,33}]
  wire  _GEN_422 = 7'h26 == reqIndex ? way1V_38 : _GEN_421; // @[ICache.scala 46:{33,33}]
  wire  _GEN_423 = 7'h27 == reqIndex ? way1V_39 : _GEN_422; // @[ICache.scala 46:{33,33}]
  wire  _GEN_424 = 7'h28 == reqIndex ? way1V_40 : _GEN_423; // @[ICache.scala 46:{33,33}]
  wire  _GEN_425 = 7'h29 == reqIndex ? way1V_41 : _GEN_424; // @[ICache.scala 46:{33,33}]
  wire  _GEN_426 = 7'h2a == reqIndex ? way1V_42 : _GEN_425; // @[ICache.scala 46:{33,33}]
  wire  _GEN_427 = 7'h2b == reqIndex ? way1V_43 : _GEN_426; // @[ICache.scala 46:{33,33}]
  wire  _GEN_428 = 7'h2c == reqIndex ? way1V_44 : _GEN_427; // @[ICache.scala 46:{33,33}]
  wire  _GEN_429 = 7'h2d == reqIndex ? way1V_45 : _GEN_428; // @[ICache.scala 46:{33,33}]
  wire  _GEN_430 = 7'h2e == reqIndex ? way1V_46 : _GEN_429; // @[ICache.scala 46:{33,33}]
  wire  _GEN_431 = 7'h2f == reqIndex ? way1V_47 : _GEN_430; // @[ICache.scala 46:{33,33}]
  wire  _GEN_432 = 7'h30 == reqIndex ? way1V_48 : _GEN_431; // @[ICache.scala 46:{33,33}]
  wire  _GEN_433 = 7'h31 == reqIndex ? way1V_49 : _GEN_432; // @[ICache.scala 46:{33,33}]
  wire  _GEN_434 = 7'h32 == reqIndex ? way1V_50 : _GEN_433; // @[ICache.scala 46:{33,33}]
  wire  _GEN_435 = 7'h33 == reqIndex ? way1V_51 : _GEN_434; // @[ICache.scala 46:{33,33}]
  wire  _GEN_436 = 7'h34 == reqIndex ? way1V_52 : _GEN_435; // @[ICache.scala 46:{33,33}]
  wire  _GEN_437 = 7'h35 == reqIndex ? way1V_53 : _GEN_436; // @[ICache.scala 46:{33,33}]
  wire  _GEN_438 = 7'h36 == reqIndex ? way1V_54 : _GEN_437; // @[ICache.scala 46:{33,33}]
  wire  _GEN_439 = 7'h37 == reqIndex ? way1V_55 : _GEN_438; // @[ICache.scala 46:{33,33}]
  wire  _GEN_440 = 7'h38 == reqIndex ? way1V_56 : _GEN_439; // @[ICache.scala 46:{33,33}]
  wire  _GEN_441 = 7'h39 == reqIndex ? way1V_57 : _GEN_440; // @[ICache.scala 46:{33,33}]
  wire  _GEN_442 = 7'h3a == reqIndex ? way1V_58 : _GEN_441; // @[ICache.scala 46:{33,33}]
  wire  _GEN_443 = 7'h3b == reqIndex ? way1V_59 : _GEN_442; // @[ICache.scala 46:{33,33}]
  wire  _GEN_444 = 7'h3c == reqIndex ? way1V_60 : _GEN_443; // @[ICache.scala 46:{33,33}]
  wire  _GEN_445 = 7'h3d == reqIndex ? way1V_61 : _GEN_444; // @[ICache.scala 46:{33,33}]
  wire  _GEN_446 = 7'h3e == reqIndex ? way1V_62 : _GEN_445; // @[ICache.scala 46:{33,33}]
  wire  _GEN_447 = 7'h3f == reqIndex ? way1V_63 : _GEN_446; // @[ICache.scala 46:{33,33}]
  wire  _GEN_448 = 7'h40 == reqIndex ? way1V_64 : _GEN_447; // @[ICache.scala 46:{33,33}]
  wire  _GEN_449 = 7'h41 == reqIndex ? way1V_65 : _GEN_448; // @[ICache.scala 46:{33,33}]
  wire  _GEN_450 = 7'h42 == reqIndex ? way1V_66 : _GEN_449; // @[ICache.scala 46:{33,33}]
  wire  _GEN_451 = 7'h43 == reqIndex ? way1V_67 : _GEN_450; // @[ICache.scala 46:{33,33}]
  wire  _GEN_452 = 7'h44 == reqIndex ? way1V_68 : _GEN_451; // @[ICache.scala 46:{33,33}]
  wire  _GEN_453 = 7'h45 == reqIndex ? way1V_69 : _GEN_452; // @[ICache.scala 46:{33,33}]
  wire  _GEN_454 = 7'h46 == reqIndex ? way1V_70 : _GEN_453; // @[ICache.scala 46:{33,33}]
  wire  _GEN_455 = 7'h47 == reqIndex ? way1V_71 : _GEN_454; // @[ICache.scala 46:{33,33}]
  wire  _GEN_456 = 7'h48 == reqIndex ? way1V_72 : _GEN_455; // @[ICache.scala 46:{33,33}]
  wire  _GEN_457 = 7'h49 == reqIndex ? way1V_73 : _GEN_456; // @[ICache.scala 46:{33,33}]
  wire  _GEN_458 = 7'h4a == reqIndex ? way1V_74 : _GEN_457; // @[ICache.scala 46:{33,33}]
  wire  _GEN_459 = 7'h4b == reqIndex ? way1V_75 : _GEN_458; // @[ICache.scala 46:{33,33}]
  wire  _GEN_460 = 7'h4c == reqIndex ? way1V_76 : _GEN_459; // @[ICache.scala 46:{33,33}]
  wire  _GEN_461 = 7'h4d == reqIndex ? way1V_77 : _GEN_460; // @[ICache.scala 46:{33,33}]
  wire  _GEN_462 = 7'h4e == reqIndex ? way1V_78 : _GEN_461; // @[ICache.scala 46:{33,33}]
  wire  _GEN_463 = 7'h4f == reqIndex ? way1V_79 : _GEN_462; // @[ICache.scala 46:{33,33}]
  wire  _GEN_464 = 7'h50 == reqIndex ? way1V_80 : _GEN_463; // @[ICache.scala 46:{33,33}]
  wire  _GEN_465 = 7'h51 == reqIndex ? way1V_81 : _GEN_464; // @[ICache.scala 46:{33,33}]
  wire  _GEN_466 = 7'h52 == reqIndex ? way1V_82 : _GEN_465; // @[ICache.scala 46:{33,33}]
  wire  _GEN_467 = 7'h53 == reqIndex ? way1V_83 : _GEN_466; // @[ICache.scala 46:{33,33}]
  wire  _GEN_468 = 7'h54 == reqIndex ? way1V_84 : _GEN_467; // @[ICache.scala 46:{33,33}]
  wire  _GEN_469 = 7'h55 == reqIndex ? way1V_85 : _GEN_468; // @[ICache.scala 46:{33,33}]
  wire  _GEN_470 = 7'h56 == reqIndex ? way1V_86 : _GEN_469; // @[ICache.scala 46:{33,33}]
  wire  _GEN_471 = 7'h57 == reqIndex ? way1V_87 : _GEN_470; // @[ICache.scala 46:{33,33}]
  wire  _GEN_472 = 7'h58 == reqIndex ? way1V_88 : _GEN_471; // @[ICache.scala 46:{33,33}]
  wire  _GEN_473 = 7'h59 == reqIndex ? way1V_89 : _GEN_472; // @[ICache.scala 46:{33,33}]
  wire  _GEN_474 = 7'h5a == reqIndex ? way1V_90 : _GEN_473; // @[ICache.scala 46:{33,33}]
  wire  _GEN_475 = 7'h5b == reqIndex ? way1V_91 : _GEN_474; // @[ICache.scala 46:{33,33}]
  wire  _GEN_476 = 7'h5c == reqIndex ? way1V_92 : _GEN_475; // @[ICache.scala 46:{33,33}]
  wire  _GEN_477 = 7'h5d == reqIndex ? way1V_93 : _GEN_476; // @[ICache.scala 46:{33,33}]
  wire  _GEN_478 = 7'h5e == reqIndex ? way1V_94 : _GEN_477; // @[ICache.scala 46:{33,33}]
  wire  _GEN_479 = 7'h5f == reqIndex ? way1V_95 : _GEN_478; // @[ICache.scala 46:{33,33}]
  wire  _GEN_480 = 7'h60 == reqIndex ? way1V_96 : _GEN_479; // @[ICache.scala 46:{33,33}]
  wire  _GEN_481 = 7'h61 == reqIndex ? way1V_97 : _GEN_480; // @[ICache.scala 46:{33,33}]
  wire  _GEN_482 = 7'h62 == reqIndex ? way1V_98 : _GEN_481; // @[ICache.scala 46:{33,33}]
  wire  _GEN_483 = 7'h63 == reqIndex ? way1V_99 : _GEN_482; // @[ICache.scala 46:{33,33}]
  wire  _GEN_484 = 7'h64 == reqIndex ? way1V_100 : _GEN_483; // @[ICache.scala 46:{33,33}]
  wire  _GEN_485 = 7'h65 == reqIndex ? way1V_101 : _GEN_484; // @[ICache.scala 46:{33,33}]
  wire  _GEN_486 = 7'h66 == reqIndex ? way1V_102 : _GEN_485; // @[ICache.scala 46:{33,33}]
  wire  _GEN_487 = 7'h67 == reqIndex ? way1V_103 : _GEN_486; // @[ICache.scala 46:{33,33}]
  wire  _GEN_488 = 7'h68 == reqIndex ? way1V_104 : _GEN_487; // @[ICache.scala 46:{33,33}]
  wire  _GEN_489 = 7'h69 == reqIndex ? way1V_105 : _GEN_488; // @[ICache.scala 46:{33,33}]
  wire  _GEN_490 = 7'h6a == reqIndex ? way1V_106 : _GEN_489; // @[ICache.scala 46:{33,33}]
  wire  _GEN_491 = 7'h6b == reqIndex ? way1V_107 : _GEN_490; // @[ICache.scala 46:{33,33}]
  wire  _GEN_492 = 7'h6c == reqIndex ? way1V_108 : _GEN_491; // @[ICache.scala 46:{33,33}]
  wire  _GEN_493 = 7'h6d == reqIndex ? way1V_109 : _GEN_492; // @[ICache.scala 46:{33,33}]
  wire  _GEN_494 = 7'h6e == reqIndex ? way1V_110 : _GEN_493; // @[ICache.scala 46:{33,33}]
  wire  _GEN_495 = 7'h6f == reqIndex ? way1V_111 : _GEN_494; // @[ICache.scala 46:{33,33}]
  wire  _GEN_496 = 7'h70 == reqIndex ? way1V_112 : _GEN_495; // @[ICache.scala 46:{33,33}]
  wire  _GEN_497 = 7'h71 == reqIndex ? way1V_113 : _GEN_496; // @[ICache.scala 46:{33,33}]
  wire  _GEN_498 = 7'h72 == reqIndex ? way1V_114 : _GEN_497; // @[ICache.scala 46:{33,33}]
  wire  _GEN_499 = 7'h73 == reqIndex ? way1V_115 : _GEN_498; // @[ICache.scala 46:{33,33}]
  wire  _GEN_500 = 7'h74 == reqIndex ? way1V_116 : _GEN_499; // @[ICache.scala 46:{33,33}]
  wire  _GEN_501 = 7'h75 == reqIndex ? way1V_117 : _GEN_500; // @[ICache.scala 46:{33,33}]
  wire  _GEN_502 = 7'h76 == reqIndex ? way1V_118 : _GEN_501; // @[ICache.scala 46:{33,33}]
  wire  _GEN_503 = 7'h77 == reqIndex ? way1V_119 : _GEN_502; // @[ICache.scala 46:{33,33}]
  wire  _GEN_504 = 7'h78 == reqIndex ? way1V_120 : _GEN_503; // @[ICache.scala 46:{33,33}]
  wire  _GEN_505 = 7'h79 == reqIndex ? way1V_121 : _GEN_504; // @[ICache.scala 46:{33,33}]
  wire  _GEN_506 = 7'h7a == reqIndex ? way1V_122 : _GEN_505; // @[ICache.scala 46:{33,33}]
  wire  _GEN_507 = 7'h7b == reqIndex ? way1V_123 : _GEN_506; // @[ICache.scala 46:{33,33}]
  wire  _GEN_508 = 7'h7c == reqIndex ? way1V_124 : _GEN_507; // @[ICache.scala 46:{33,33}]
  wire  _GEN_509 = 7'h7d == reqIndex ? way1V_125 : _GEN_508; // @[ICache.scala 46:{33,33}]
  wire  _GEN_510 = 7'h7e == reqIndex ? way1V_126 : _GEN_509; // @[ICache.scala 46:{33,33}]
  wire  _GEN_511 = 7'h7f == reqIndex ? way1V_127 : _GEN_510; // @[ICache.scala 46:{33,33}]
  wire  way1Hit = _GEN_511 & _GEN_383 == reqTag; // @[ICache.scala 46:33]
  wire [7:0] _cacheRIndex_T = {1'h0,reqIndex}; // @[Cat.scala 31:58]
  wire [7:0] _cacheRIndex_T_1 = {1'h1,reqIndex}; // @[Cat.scala 31:58]
  wire [7:0] cacheRIndex = way0Hit ? _cacheRIndex_T : _cacheRIndex_T_1; // @[ICache.scala 47:24]
  wire  cacheHitEn = way0Hit | way1Hit; // @[ICache.scala 49:28]
  wire  sFillEn = state == 2'h3; // @[ICache.scala 104:23]
  wire  _GEN_520 = 7'h1 == reqIndex ? way0Age_1 : way0Age_0; // @[ICache.scala 106:{38,38}]
  wire  _GEN_521 = 7'h2 == reqIndex ? way0Age_2 : _GEN_520; // @[ICache.scala 106:{38,38}]
  wire  _GEN_522 = 7'h3 == reqIndex ? way0Age_3 : _GEN_521; // @[ICache.scala 106:{38,38}]
  wire  _GEN_523 = 7'h4 == reqIndex ? way0Age_4 : _GEN_522; // @[ICache.scala 106:{38,38}]
  wire  _GEN_524 = 7'h5 == reqIndex ? way0Age_5 : _GEN_523; // @[ICache.scala 106:{38,38}]
  wire  _GEN_525 = 7'h6 == reqIndex ? way0Age_6 : _GEN_524; // @[ICache.scala 106:{38,38}]
  wire  _GEN_526 = 7'h7 == reqIndex ? way0Age_7 : _GEN_525; // @[ICache.scala 106:{38,38}]
  wire  _GEN_527 = 7'h8 == reqIndex ? way0Age_8 : _GEN_526; // @[ICache.scala 106:{38,38}]
  wire  _GEN_528 = 7'h9 == reqIndex ? way0Age_9 : _GEN_527; // @[ICache.scala 106:{38,38}]
  wire  _GEN_529 = 7'ha == reqIndex ? way0Age_10 : _GEN_528; // @[ICache.scala 106:{38,38}]
  wire  _GEN_530 = 7'hb == reqIndex ? way0Age_11 : _GEN_529; // @[ICache.scala 106:{38,38}]
  wire  _GEN_531 = 7'hc == reqIndex ? way0Age_12 : _GEN_530; // @[ICache.scala 106:{38,38}]
  wire  _GEN_532 = 7'hd == reqIndex ? way0Age_13 : _GEN_531; // @[ICache.scala 106:{38,38}]
  wire  _GEN_533 = 7'he == reqIndex ? way0Age_14 : _GEN_532; // @[ICache.scala 106:{38,38}]
  wire  _GEN_534 = 7'hf == reqIndex ? way0Age_15 : _GEN_533; // @[ICache.scala 106:{38,38}]
  wire  _GEN_535 = 7'h10 == reqIndex ? way0Age_16 : _GEN_534; // @[ICache.scala 106:{38,38}]
  wire  _GEN_536 = 7'h11 == reqIndex ? way0Age_17 : _GEN_535; // @[ICache.scala 106:{38,38}]
  wire  _GEN_537 = 7'h12 == reqIndex ? way0Age_18 : _GEN_536; // @[ICache.scala 106:{38,38}]
  wire  _GEN_538 = 7'h13 == reqIndex ? way0Age_19 : _GEN_537; // @[ICache.scala 106:{38,38}]
  wire  _GEN_539 = 7'h14 == reqIndex ? way0Age_20 : _GEN_538; // @[ICache.scala 106:{38,38}]
  wire  _GEN_540 = 7'h15 == reqIndex ? way0Age_21 : _GEN_539; // @[ICache.scala 106:{38,38}]
  wire  _GEN_541 = 7'h16 == reqIndex ? way0Age_22 : _GEN_540; // @[ICache.scala 106:{38,38}]
  wire  _GEN_542 = 7'h17 == reqIndex ? way0Age_23 : _GEN_541; // @[ICache.scala 106:{38,38}]
  wire  _GEN_543 = 7'h18 == reqIndex ? way0Age_24 : _GEN_542; // @[ICache.scala 106:{38,38}]
  wire  _GEN_544 = 7'h19 == reqIndex ? way0Age_25 : _GEN_543; // @[ICache.scala 106:{38,38}]
  wire  _GEN_545 = 7'h1a == reqIndex ? way0Age_26 : _GEN_544; // @[ICache.scala 106:{38,38}]
  wire  _GEN_546 = 7'h1b == reqIndex ? way0Age_27 : _GEN_545; // @[ICache.scala 106:{38,38}]
  wire  _GEN_547 = 7'h1c == reqIndex ? way0Age_28 : _GEN_546; // @[ICache.scala 106:{38,38}]
  wire  _GEN_548 = 7'h1d == reqIndex ? way0Age_29 : _GEN_547; // @[ICache.scala 106:{38,38}]
  wire  _GEN_549 = 7'h1e == reqIndex ? way0Age_30 : _GEN_548; // @[ICache.scala 106:{38,38}]
  wire  _GEN_550 = 7'h1f == reqIndex ? way0Age_31 : _GEN_549; // @[ICache.scala 106:{38,38}]
  wire  _GEN_551 = 7'h20 == reqIndex ? way0Age_32 : _GEN_550; // @[ICache.scala 106:{38,38}]
  wire  _GEN_552 = 7'h21 == reqIndex ? way0Age_33 : _GEN_551; // @[ICache.scala 106:{38,38}]
  wire  _GEN_553 = 7'h22 == reqIndex ? way0Age_34 : _GEN_552; // @[ICache.scala 106:{38,38}]
  wire  _GEN_554 = 7'h23 == reqIndex ? way0Age_35 : _GEN_553; // @[ICache.scala 106:{38,38}]
  wire  _GEN_555 = 7'h24 == reqIndex ? way0Age_36 : _GEN_554; // @[ICache.scala 106:{38,38}]
  wire  _GEN_556 = 7'h25 == reqIndex ? way0Age_37 : _GEN_555; // @[ICache.scala 106:{38,38}]
  wire  _GEN_557 = 7'h26 == reqIndex ? way0Age_38 : _GEN_556; // @[ICache.scala 106:{38,38}]
  wire  _GEN_558 = 7'h27 == reqIndex ? way0Age_39 : _GEN_557; // @[ICache.scala 106:{38,38}]
  wire  _GEN_559 = 7'h28 == reqIndex ? way0Age_40 : _GEN_558; // @[ICache.scala 106:{38,38}]
  wire  _GEN_560 = 7'h29 == reqIndex ? way0Age_41 : _GEN_559; // @[ICache.scala 106:{38,38}]
  wire  _GEN_561 = 7'h2a == reqIndex ? way0Age_42 : _GEN_560; // @[ICache.scala 106:{38,38}]
  wire  _GEN_562 = 7'h2b == reqIndex ? way0Age_43 : _GEN_561; // @[ICache.scala 106:{38,38}]
  wire  _GEN_563 = 7'h2c == reqIndex ? way0Age_44 : _GEN_562; // @[ICache.scala 106:{38,38}]
  wire  _GEN_564 = 7'h2d == reqIndex ? way0Age_45 : _GEN_563; // @[ICache.scala 106:{38,38}]
  wire  _GEN_565 = 7'h2e == reqIndex ? way0Age_46 : _GEN_564; // @[ICache.scala 106:{38,38}]
  wire  _GEN_566 = 7'h2f == reqIndex ? way0Age_47 : _GEN_565; // @[ICache.scala 106:{38,38}]
  wire  _GEN_567 = 7'h30 == reqIndex ? way0Age_48 : _GEN_566; // @[ICache.scala 106:{38,38}]
  wire  _GEN_568 = 7'h31 == reqIndex ? way0Age_49 : _GEN_567; // @[ICache.scala 106:{38,38}]
  wire  _GEN_569 = 7'h32 == reqIndex ? way0Age_50 : _GEN_568; // @[ICache.scala 106:{38,38}]
  wire  _GEN_570 = 7'h33 == reqIndex ? way0Age_51 : _GEN_569; // @[ICache.scala 106:{38,38}]
  wire  _GEN_571 = 7'h34 == reqIndex ? way0Age_52 : _GEN_570; // @[ICache.scala 106:{38,38}]
  wire  _GEN_572 = 7'h35 == reqIndex ? way0Age_53 : _GEN_571; // @[ICache.scala 106:{38,38}]
  wire  _GEN_573 = 7'h36 == reqIndex ? way0Age_54 : _GEN_572; // @[ICache.scala 106:{38,38}]
  wire  _GEN_574 = 7'h37 == reqIndex ? way0Age_55 : _GEN_573; // @[ICache.scala 106:{38,38}]
  wire  _GEN_575 = 7'h38 == reqIndex ? way0Age_56 : _GEN_574; // @[ICache.scala 106:{38,38}]
  wire  _GEN_576 = 7'h39 == reqIndex ? way0Age_57 : _GEN_575; // @[ICache.scala 106:{38,38}]
  wire  _GEN_577 = 7'h3a == reqIndex ? way0Age_58 : _GEN_576; // @[ICache.scala 106:{38,38}]
  wire  _GEN_578 = 7'h3b == reqIndex ? way0Age_59 : _GEN_577; // @[ICache.scala 106:{38,38}]
  wire  _GEN_579 = 7'h3c == reqIndex ? way0Age_60 : _GEN_578; // @[ICache.scala 106:{38,38}]
  wire  _GEN_580 = 7'h3d == reqIndex ? way0Age_61 : _GEN_579; // @[ICache.scala 106:{38,38}]
  wire  _GEN_581 = 7'h3e == reqIndex ? way0Age_62 : _GEN_580; // @[ICache.scala 106:{38,38}]
  wire  _GEN_582 = 7'h3f == reqIndex ? way0Age_63 : _GEN_581; // @[ICache.scala 106:{38,38}]
  wire  _GEN_583 = 7'h40 == reqIndex ? way0Age_64 : _GEN_582; // @[ICache.scala 106:{38,38}]
  wire  _GEN_584 = 7'h41 == reqIndex ? way0Age_65 : _GEN_583; // @[ICache.scala 106:{38,38}]
  wire  _GEN_585 = 7'h42 == reqIndex ? way0Age_66 : _GEN_584; // @[ICache.scala 106:{38,38}]
  wire  _GEN_586 = 7'h43 == reqIndex ? way0Age_67 : _GEN_585; // @[ICache.scala 106:{38,38}]
  wire  _GEN_587 = 7'h44 == reqIndex ? way0Age_68 : _GEN_586; // @[ICache.scala 106:{38,38}]
  wire  _GEN_588 = 7'h45 == reqIndex ? way0Age_69 : _GEN_587; // @[ICache.scala 106:{38,38}]
  wire  _GEN_589 = 7'h46 == reqIndex ? way0Age_70 : _GEN_588; // @[ICache.scala 106:{38,38}]
  wire  _GEN_590 = 7'h47 == reqIndex ? way0Age_71 : _GEN_589; // @[ICache.scala 106:{38,38}]
  wire  _GEN_591 = 7'h48 == reqIndex ? way0Age_72 : _GEN_590; // @[ICache.scala 106:{38,38}]
  wire  _GEN_592 = 7'h49 == reqIndex ? way0Age_73 : _GEN_591; // @[ICache.scala 106:{38,38}]
  wire  _GEN_593 = 7'h4a == reqIndex ? way0Age_74 : _GEN_592; // @[ICache.scala 106:{38,38}]
  wire  _GEN_594 = 7'h4b == reqIndex ? way0Age_75 : _GEN_593; // @[ICache.scala 106:{38,38}]
  wire  _GEN_595 = 7'h4c == reqIndex ? way0Age_76 : _GEN_594; // @[ICache.scala 106:{38,38}]
  wire  _GEN_596 = 7'h4d == reqIndex ? way0Age_77 : _GEN_595; // @[ICache.scala 106:{38,38}]
  wire  _GEN_597 = 7'h4e == reqIndex ? way0Age_78 : _GEN_596; // @[ICache.scala 106:{38,38}]
  wire  _GEN_598 = 7'h4f == reqIndex ? way0Age_79 : _GEN_597; // @[ICache.scala 106:{38,38}]
  wire  _GEN_599 = 7'h50 == reqIndex ? way0Age_80 : _GEN_598; // @[ICache.scala 106:{38,38}]
  wire  _GEN_600 = 7'h51 == reqIndex ? way0Age_81 : _GEN_599; // @[ICache.scala 106:{38,38}]
  wire  _GEN_601 = 7'h52 == reqIndex ? way0Age_82 : _GEN_600; // @[ICache.scala 106:{38,38}]
  wire  _GEN_602 = 7'h53 == reqIndex ? way0Age_83 : _GEN_601; // @[ICache.scala 106:{38,38}]
  wire  _GEN_603 = 7'h54 == reqIndex ? way0Age_84 : _GEN_602; // @[ICache.scala 106:{38,38}]
  wire  _GEN_604 = 7'h55 == reqIndex ? way0Age_85 : _GEN_603; // @[ICache.scala 106:{38,38}]
  wire  _GEN_605 = 7'h56 == reqIndex ? way0Age_86 : _GEN_604; // @[ICache.scala 106:{38,38}]
  wire  _GEN_606 = 7'h57 == reqIndex ? way0Age_87 : _GEN_605; // @[ICache.scala 106:{38,38}]
  wire  _GEN_607 = 7'h58 == reqIndex ? way0Age_88 : _GEN_606; // @[ICache.scala 106:{38,38}]
  wire  _GEN_608 = 7'h59 == reqIndex ? way0Age_89 : _GEN_607; // @[ICache.scala 106:{38,38}]
  wire  _GEN_609 = 7'h5a == reqIndex ? way0Age_90 : _GEN_608; // @[ICache.scala 106:{38,38}]
  wire  _GEN_610 = 7'h5b == reqIndex ? way0Age_91 : _GEN_609; // @[ICache.scala 106:{38,38}]
  wire  _GEN_611 = 7'h5c == reqIndex ? way0Age_92 : _GEN_610; // @[ICache.scala 106:{38,38}]
  wire  _GEN_612 = 7'h5d == reqIndex ? way0Age_93 : _GEN_611; // @[ICache.scala 106:{38,38}]
  wire  _GEN_613 = 7'h5e == reqIndex ? way0Age_94 : _GEN_612; // @[ICache.scala 106:{38,38}]
  wire  _GEN_614 = 7'h5f == reqIndex ? way0Age_95 : _GEN_613; // @[ICache.scala 106:{38,38}]
  wire  _GEN_615 = 7'h60 == reqIndex ? way0Age_96 : _GEN_614; // @[ICache.scala 106:{38,38}]
  wire  _GEN_616 = 7'h61 == reqIndex ? way0Age_97 : _GEN_615; // @[ICache.scala 106:{38,38}]
  wire  _GEN_617 = 7'h62 == reqIndex ? way0Age_98 : _GEN_616; // @[ICache.scala 106:{38,38}]
  wire  _GEN_618 = 7'h63 == reqIndex ? way0Age_99 : _GEN_617; // @[ICache.scala 106:{38,38}]
  wire  _GEN_619 = 7'h64 == reqIndex ? way0Age_100 : _GEN_618; // @[ICache.scala 106:{38,38}]
  wire  _GEN_620 = 7'h65 == reqIndex ? way0Age_101 : _GEN_619; // @[ICache.scala 106:{38,38}]
  wire  _GEN_621 = 7'h66 == reqIndex ? way0Age_102 : _GEN_620; // @[ICache.scala 106:{38,38}]
  wire  _GEN_622 = 7'h67 == reqIndex ? way0Age_103 : _GEN_621; // @[ICache.scala 106:{38,38}]
  wire  _GEN_623 = 7'h68 == reqIndex ? way0Age_104 : _GEN_622; // @[ICache.scala 106:{38,38}]
  wire  _GEN_624 = 7'h69 == reqIndex ? way0Age_105 : _GEN_623; // @[ICache.scala 106:{38,38}]
  wire  _GEN_625 = 7'h6a == reqIndex ? way0Age_106 : _GEN_624; // @[ICache.scala 106:{38,38}]
  wire  _GEN_626 = 7'h6b == reqIndex ? way0Age_107 : _GEN_625; // @[ICache.scala 106:{38,38}]
  wire  _GEN_627 = 7'h6c == reqIndex ? way0Age_108 : _GEN_626; // @[ICache.scala 106:{38,38}]
  wire  _GEN_628 = 7'h6d == reqIndex ? way0Age_109 : _GEN_627; // @[ICache.scala 106:{38,38}]
  wire  _GEN_629 = 7'h6e == reqIndex ? way0Age_110 : _GEN_628; // @[ICache.scala 106:{38,38}]
  wire  _GEN_630 = 7'h6f == reqIndex ? way0Age_111 : _GEN_629; // @[ICache.scala 106:{38,38}]
  wire  _GEN_631 = 7'h70 == reqIndex ? way0Age_112 : _GEN_630; // @[ICache.scala 106:{38,38}]
  wire  _GEN_632 = 7'h71 == reqIndex ? way0Age_113 : _GEN_631; // @[ICache.scala 106:{38,38}]
  wire  _GEN_633 = 7'h72 == reqIndex ? way0Age_114 : _GEN_632; // @[ICache.scala 106:{38,38}]
  wire  _GEN_634 = 7'h73 == reqIndex ? way0Age_115 : _GEN_633; // @[ICache.scala 106:{38,38}]
  wire  _GEN_635 = 7'h74 == reqIndex ? way0Age_116 : _GEN_634; // @[ICache.scala 106:{38,38}]
  wire  _GEN_636 = 7'h75 == reqIndex ? way0Age_117 : _GEN_635; // @[ICache.scala 106:{38,38}]
  wire  _GEN_637 = 7'h76 == reqIndex ? way0Age_118 : _GEN_636; // @[ICache.scala 106:{38,38}]
  wire  _GEN_638 = 7'h77 == reqIndex ? way0Age_119 : _GEN_637; // @[ICache.scala 106:{38,38}]
  wire  _GEN_639 = 7'h78 == reqIndex ? way0Age_120 : _GEN_638; // @[ICache.scala 106:{38,38}]
  wire  _GEN_640 = 7'h79 == reqIndex ? way0Age_121 : _GEN_639; // @[ICache.scala 106:{38,38}]
  wire  _GEN_641 = 7'h7a == reqIndex ? way0Age_122 : _GEN_640; // @[ICache.scala 106:{38,38}]
  wire  _GEN_642 = 7'h7b == reqIndex ? way0Age_123 : _GEN_641; // @[ICache.scala 106:{38,38}]
  wire  _GEN_643 = 7'h7c == reqIndex ? way0Age_124 : _GEN_642; // @[ICache.scala 106:{38,38}]
  wire  _GEN_644 = 7'h7d == reqIndex ? way0Age_125 : _GEN_643; // @[ICache.scala 106:{38,38}]
  wire  _GEN_645 = 7'h7e == reqIndex ? way0Age_126 : _GEN_644; // @[ICache.scala 106:{38,38}]
  wire  _GEN_646 = 7'h7f == reqIndex ? way0Age_127 : _GEN_645; // @[ICache.scala 106:{38,38}]
  wire  ageWay0En = ~_GEN_646 & sFillEn; // @[ICache.scala 106:47]
  wire  cacheLineWay = ageWay0En ? 1'h0 : 1'h1; // @[ICache.scala 108:25]
  wire [7:0] cacheWIndex = {cacheLineWay,reqIndex}; // @[Cat.scala 31:58]
  wire [1:0] _GEN_514 = io_out_inst_ready ? 2'h3 : state; // @[ICache.scala 76:28 77:15 38:22]
  wire [1:0] _GEN_515 = 2'h3 == state ? 2'h1 : state; // @[ICache.scala 60:17 82:15 38:22]
  wire  sReadEn = state == 2'h1; // @[ICache.scala 86:23]
  wire [127:0] cacheRData = req_Q;
  wire [127:0] rData = sReadEn & cacheHitEn ? cacheRData : 128'h0; // @[ICache.scala 87:18]
  wire [31:0] _io_imem_inst_read_T_6 = 2'h1 == reqOff[3:2] ? rData[63:32] : rData[31:0]; // @[Mux.scala 81:58]
  wire [31:0] _io_imem_inst_read_T_8 = 2'h2 == reqOff[3:2] ? rData[95:64] : _io_imem_inst_read_T_6; // @[Mux.scala 81:58]
  wire  sAxiEn = state == 2'h2; // @[ICache.scala 96:22]
  wire  _GEN_648 = 7'h1 == reqIndex ? way1Age_1 : way1Age_0; // @[ICache.scala 107:{38,38}]
  wire  _GEN_649 = 7'h2 == reqIndex ? way1Age_2 : _GEN_648; // @[ICache.scala 107:{38,38}]
  wire  _GEN_650 = 7'h3 == reqIndex ? way1Age_3 : _GEN_649; // @[ICache.scala 107:{38,38}]
  wire  _GEN_651 = 7'h4 == reqIndex ? way1Age_4 : _GEN_650; // @[ICache.scala 107:{38,38}]
  wire  _GEN_652 = 7'h5 == reqIndex ? way1Age_5 : _GEN_651; // @[ICache.scala 107:{38,38}]
  wire  _GEN_653 = 7'h6 == reqIndex ? way1Age_6 : _GEN_652; // @[ICache.scala 107:{38,38}]
  wire  _GEN_654 = 7'h7 == reqIndex ? way1Age_7 : _GEN_653; // @[ICache.scala 107:{38,38}]
  wire  _GEN_655 = 7'h8 == reqIndex ? way1Age_8 : _GEN_654; // @[ICache.scala 107:{38,38}]
  wire  _GEN_656 = 7'h9 == reqIndex ? way1Age_9 : _GEN_655; // @[ICache.scala 107:{38,38}]
  wire  _GEN_657 = 7'ha == reqIndex ? way1Age_10 : _GEN_656; // @[ICache.scala 107:{38,38}]
  wire  _GEN_658 = 7'hb == reqIndex ? way1Age_11 : _GEN_657; // @[ICache.scala 107:{38,38}]
  wire  _GEN_659 = 7'hc == reqIndex ? way1Age_12 : _GEN_658; // @[ICache.scala 107:{38,38}]
  wire  _GEN_660 = 7'hd == reqIndex ? way1Age_13 : _GEN_659; // @[ICache.scala 107:{38,38}]
  wire  _GEN_661 = 7'he == reqIndex ? way1Age_14 : _GEN_660; // @[ICache.scala 107:{38,38}]
  wire  _GEN_662 = 7'hf == reqIndex ? way1Age_15 : _GEN_661; // @[ICache.scala 107:{38,38}]
  wire  _GEN_663 = 7'h10 == reqIndex ? way1Age_16 : _GEN_662; // @[ICache.scala 107:{38,38}]
  wire  _GEN_664 = 7'h11 == reqIndex ? way1Age_17 : _GEN_663; // @[ICache.scala 107:{38,38}]
  wire  _GEN_665 = 7'h12 == reqIndex ? way1Age_18 : _GEN_664; // @[ICache.scala 107:{38,38}]
  wire  _GEN_666 = 7'h13 == reqIndex ? way1Age_19 : _GEN_665; // @[ICache.scala 107:{38,38}]
  wire  _GEN_667 = 7'h14 == reqIndex ? way1Age_20 : _GEN_666; // @[ICache.scala 107:{38,38}]
  wire  _GEN_668 = 7'h15 == reqIndex ? way1Age_21 : _GEN_667; // @[ICache.scala 107:{38,38}]
  wire  _GEN_669 = 7'h16 == reqIndex ? way1Age_22 : _GEN_668; // @[ICache.scala 107:{38,38}]
  wire  _GEN_670 = 7'h17 == reqIndex ? way1Age_23 : _GEN_669; // @[ICache.scala 107:{38,38}]
  wire  _GEN_671 = 7'h18 == reqIndex ? way1Age_24 : _GEN_670; // @[ICache.scala 107:{38,38}]
  wire  _GEN_672 = 7'h19 == reqIndex ? way1Age_25 : _GEN_671; // @[ICache.scala 107:{38,38}]
  wire  _GEN_673 = 7'h1a == reqIndex ? way1Age_26 : _GEN_672; // @[ICache.scala 107:{38,38}]
  wire  _GEN_674 = 7'h1b == reqIndex ? way1Age_27 : _GEN_673; // @[ICache.scala 107:{38,38}]
  wire  _GEN_675 = 7'h1c == reqIndex ? way1Age_28 : _GEN_674; // @[ICache.scala 107:{38,38}]
  wire  _GEN_676 = 7'h1d == reqIndex ? way1Age_29 : _GEN_675; // @[ICache.scala 107:{38,38}]
  wire  _GEN_677 = 7'h1e == reqIndex ? way1Age_30 : _GEN_676; // @[ICache.scala 107:{38,38}]
  wire  _GEN_678 = 7'h1f == reqIndex ? way1Age_31 : _GEN_677; // @[ICache.scala 107:{38,38}]
  wire  _GEN_679 = 7'h20 == reqIndex ? way1Age_32 : _GEN_678; // @[ICache.scala 107:{38,38}]
  wire  _GEN_680 = 7'h21 == reqIndex ? way1Age_33 : _GEN_679; // @[ICache.scala 107:{38,38}]
  wire  _GEN_681 = 7'h22 == reqIndex ? way1Age_34 : _GEN_680; // @[ICache.scala 107:{38,38}]
  wire  _GEN_682 = 7'h23 == reqIndex ? way1Age_35 : _GEN_681; // @[ICache.scala 107:{38,38}]
  wire  _GEN_683 = 7'h24 == reqIndex ? way1Age_36 : _GEN_682; // @[ICache.scala 107:{38,38}]
  wire  _GEN_684 = 7'h25 == reqIndex ? way1Age_37 : _GEN_683; // @[ICache.scala 107:{38,38}]
  wire  _GEN_685 = 7'h26 == reqIndex ? way1Age_38 : _GEN_684; // @[ICache.scala 107:{38,38}]
  wire  _GEN_686 = 7'h27 == reqIndex ? way1Age_39 : _GEN_685; // @[ICache.scala 107:{38,38}]
  wire  _GEN_687 = 7'h28 == reqIndex ? way1Age_40 : _GEN_686; // @[ICache.scala 107:{38,38}]
  wire  _GEN_688 = 7'h29 == reqIndex ? way1Age_41 : _GEN_687; // @[ICache.scala 107:{38,38}]
  wire  _GEN_689 = 7'h2a == reqIndex ? way1Age_42 : _GEN_688; // @[ICache.scala 107:{38,38}]
  wire  _GEN_690 = 7'h2b == reqIndex ? way1Age_43 : _GEN_689; // @[ICache.scala 107:{38,38}]
  wire  _GEN_691 = 7'h2c == reqIndex ? way1Age_44 : _GEN_690; // @[ICache.scala 107:{38,38}]
  wire  _GEN_692 = 7'h2d == reqIndex ? way1Age_45 : _GEN_691; // @[ICache.scala 107:{38,38}]
  wire  _GEN_693 = 7'h2e == reqIndex ? way1Age_46 : _GEN_692; // @[ICache.scala 107:{38,38}]
  wire  _GEN_694 = 7'h2f == reqIndex ? way1Age_47 : _GEN_693; // @[ICache.scala 107:{38,38}]
  wire  _GEN_695 = 7'h30 == reqIndex ? way1Age_48 : _GEN_694; // @[ICache.scala 107:{38,38}]
  wire  _GEN_696 = 7'h31 == reqIndex ? way1Age_49 : _GEN_695; // @[ICache.scala 107:{38,38}]
  wire  _GEN_697 = 7'h32 == reqIndex ? way1Age_50 : _GEN_696; // @[ICache.scala 107:{38,38}]
  wire  _GEN_698 = 7'h33 == reqIndex ? way1Age_51 : _GEN_697; // @[ICache.scala 107:{38,38}]
  wire  _GEN_699 = 7'h34 == reqIndex ? way1Age_52 : _GEN_698; // @[ICache.scala 107:{38,38}]
  wire  _GEN_700 = 7'h35 == reqIndex ? way1Age_53 : _GEN_699; // @[ICache.scala 107:{38,38}]
  wire  _GEN_701 = 7'h36 == reqIndex ? way1Age_54 : _GEN_700; // @[ICache.scala 107:{38,38}]
  wire  _GEN_702 = 7'h37 == reqIndex ? way1Age_55 : _GEN_701; // @[ICache.scala 107:{38,38}]
  wire  _GEN_703 = 7'h38 == reqIndex ? way1Age_56 : _GEN_702; // @[ICache.scala 107:{38,38}]
  wire  _GEN_704 = 7'h39 == reqIndex ? way1Age_57 : _GEN_703; // @[ICache.scala 107:{38,38}]
  wire  _GEN_705 = 7'h3a == reqIndex ? way1Age_58 : _GEN_704; // @[ICache.scala 107:{38,38}]
  wire  _GEN_706 = 7'h3b == reqIndex ? way1Age_59 : _GEN_705; // @[ICache.scala 107:{38,38}]
  wire  _GEN_707 = 7'h3c == reqIndex ? way1Age_60 : _GEN_706; // @[ICache.scala 107:{38,38}]
  wire  _GEN_708 = 7'h3d == reqIndex ? way1Age_61 : _GEN_707; // @[ICache.scala 107:{38,38}]
  wire  _GEN_709 = 7'h3e == reqIndex ? way1Age_62 : _GEN_708; // @[ICache.scala 107:{38,38}]
  wire  _GEN_710 = 7'h3f == reqIndex ? way1Age_63 : _GEN_709; // @[ICache.scala 107:{38,38}]
  wire  _GEN_711 = 7'h40 == reqIndex ? way1Age_64 : _GEN_710; // @[ICache.scala 107:{38,38}]
  wire  _GEN_712 = 7'h41 == reqIndex ? way1Age_65 : _GEN_711; // @[ICache.scala 107:{38,38}]
  wire  _GEN_713 = 7'h42 == reqIndex ? way1Age_66 : _GEN_712; // @[ICache.scala 107:{38,38}]
  wire  _GEN_714 = 7'h43 == reqIndex ? way1Age_67 : _GEN_713; // @[ICache.scala 107:{38,38}]
  wire  _GEN_715 = 7'h44 == reqIndex ? way1Age_68 : _GEN_714; // @[ICache.scala 107:{38,38}]
  wire  _GEN_716 = 7'h45 == reqIndex ? way1Age_69 : _GEN_715; // @[ICache.scala 107:{38,38}]
  wire  _GEN_717 = 7'h46 == reqIndex ? way1Age_70 : _GEN_716; // @[ICache.scala 107:{38,38}]
  wire  _GEN_718 = 7'h47 == reqIndex ? way1Age_71 : _GEN_717; // @[ICache.scala 107:{38,38}]
  wire  _GEN_719 = 7'h48 == reqIndex ? way1Age_72 : _GEN_718; // @[ICache.scala 107:{38,38}]
  wire  _GEN_720 = 7'h49 == reqIndex ? way1Age_73 : _GEN_719; // @[ICache.scala 107:{38,38}]
  wire  _GEN_721 = 7'h4a == reqIndex ? way1Age_74 : _GEN_720; // @[ICache.scala 107:{38,38}]
  wire  _GEN_722 = 7'h4b == reqIndex ? way1Age_75 : _GEN_721; // @[ICache.scala 107:{38,38}]
  wire  _GEN_723 = 7'h4c == reqIndex ? way1Age_76 : _GEN_722; // @[ICache.scala 107:{38,38}]
  wire  _GEN_724 = 7'h4d == reqIndex ? way1Age_77 : _GEN_723; // @[ICache.scala 107:{38,38}]
  wire  _GEN_725 = 7'h4e == reqIndex ? way1Age_78 : _GEN_724; // @[ICache.scala 107:{38,38}]
  wire  _GEN_726 = 7'h4f == reqIndex ? way1Age_79 : _GEN_725; // @[ICache.scala 107:{38,38}]
  wire  _GEN_727 = 7'h50 == reqIndex ? way1Age_80 : _GEN_726; // @[ICache.scala 107:{38,38}]
  wire  _GEN_728 = 7'h51 == reqIndex ? way1Age_81 : _GEN_727; // @[ICache.scala 107:{38,38}]
  wire  _GEN_729 = 7'h52 == reqIndex ? way1Age_82 : _GEN_728; // @[ICache.scala 107:{38,38}]
  wire  _GEN_730 = 7'h53 == reqIndex ? way1Age_83 : _GEN_729; // @[ICache.scala 107:{38,38}]
  wire  _GEN_731 = 7'h54 == reqIndex ? way1Age_84 : _GEN_730; // @[ICache.scala 107:{38,38}]
  wire  _GEN_732 = 7'h55 == reqIndex ? way1Age_85 : _GEN_731; // @[ICache.scala 107:{38,38}]
  wire  _GEN_733 = 7'h56 == reqIndex ? way1Age_86 : _GEN_732; // @[ICache.scala 107:{38,38}]
  wire  _GEN_734 = 7'h57 == reqIndex ? way1Age_87 : _GEN_733; // @[ICache.scala 107:{38,38}]
  wire  _GEN_735 = 7'h58 == reqIndex ? way1Age_88 : _GEN_734; // @[ICache.scala 107:{38,38}]
  wire  _GEN_736 = 7'h59 == reqIndex ? way1Age_89 : _GEN_735; // @[ICache.scala 107:{38,38}]
  wire  _GEN_737 = 7'h5a == reqIndex ? way1Age_90 : _GEN_736; // @[ICache.scala 107:{38,38}]
  wire  _GEN_738 = 7'h5b == reqIndex ? way1Age_91 : _GEN_737; // @[ICache.scala 107:{38,38}]
  wire  _GEN_739 = 7'h5c == reqIndex ? way1Age_92 : _GEN_738; // @[ICache.scala 107:{38,38}]
  wire  _GEN_740 = 7'h5d == reqIndex ? way1Age_93 : _GEN_739; // @[ICache.scala 107:{38,38}]
  wire  _GEN_741 = 7'h5e == reqIndex ? way1Age_94 : _GEN_740; // @[ICache.scala 107:{38,38}]
  wire  _GEN_742 = 7'h5f == reqIndex ? way1Age_95 : _GEN_741; // @[ICache.scala 107:{38,38}]
  wire  _GEN_743 = 7'h60 == reqIndex ? way1Age_96 : _GEN_742; // @[ICache.scala 107:{38,38}]
  wire  _GEN_744 = 7'h61 == reqIndex ? way1Age_97 : _GEN_743; // @[ICache.scala 107:{38,38}]
  wire  _GEN_745 = 7'h62 == reqIndex ? way1Age_98 : _GEN_744; // @[ICache.scala 107:{38,38}]
  wire  _GEN_746 = 7'h63 == reqIndex ? way1Age_99 : _GEN_745; // @[ICache.scala 107:{38,38}]
  wire  _GEN_747 = 7'h64 == reqIndex ? way1Age_100 : _GEN_746; // @[ICache.scala 107:{38,38}]
  wire  _GEN_748 = 7'h65 == reqIndex ? way1Age_101 : _GEN_747; // @[ICache.scala 107:{38,38}]
  wire  _GEN_749 = 7'h66 == reqIndex ? way1Age_102 : _GEN_748; // @[ICache.scala 107:{38,38}]
  wire  _GEN_750 = 7'h67 == reqIndex ? way1Age_103 : _GEN_749; // @[ICache.scala 107:{38,38}]
  wire  _GEN_751 = 7'h68 == reqIndex ? way1Age_104 : _GEN_750; // @[ICache.scala 107:{38,38}]
  wire  _GEN_752 = 7'h69 == reqIndex ? way1Age_105 : _GEN_751; // @[ICache.scala 107:{38,38}]
  wire  _GEN_753 = 7'h6a == reqIndex ? way1Age_106 : _GEN_752; // @[ICache.scala 107:{38,38}]
  wire  _GEN_754 = 7'h6b == reqIndex ? way1Age_107 : _GEN_753; // @[ICache.scala 107:{38,38}]
  wire  _GEN_755 = 7'h6c == reqIndex ? way1Age_108 : _GEN_754; // @[ICache.scala 107:{38,38}]
  wire  _GEN_756 = 7'h6d == reqIndex ? way1Age_109 : _GEN_755; // @[ICache.scala 107:{38,38}]
  wire  _GEN_757 = 7'h6e == reqIndex ? way1Age_110 : _GEN_756; // @[ICache.scala 107:{38,38}]
  wire  _GEN_758 = 7'h6f == reqIndex ? way1Age_111 : _GEN_757; // @[ICache.scala 107:{38,38}]
  wire  _GEN_759 = 7'h70 == reqIndex ? way1Age_112 : _GEN_758; // @[ICache.scala 107:{38,38}]
  wire  _GEN_760 = 7'h71 == reqIndex ? way1Age_113 : _GEN_759; // @[ICache.scala 107:{38,38}]
  wire  _GEN_761 = 7'h72 == reqIndex ? way1Age_114 : _GEN_760; // @[ICache.scala 107:{38,38}]
  wire  _GEN_762 = 7'h73 == reqIndex ? way1Age_115 : _GEN_761; // @[ICache.scala 107:{38,38}]
  wire  _GEN_763 = 7'h74 == reqIndex ? way1Age_116 : _GEN_762; // @[ICache.scala 107:{38,38}]
  wire  _GEN_764 = 7'h75 == reqIndex ? way1Age_117 : _GEN_763; // @[ICache.scala 107:{38,38}]
  wire  _GEN_765 = 7'h76 == reqIndex ? way1Age_118 : _GEN_764; // @[ICache.scala 107:{38,38}]
  wire  _GEN_766 = 7'h77 == reqIndex ? way1Age_119 : _GEN_765; // @[ICache.scala 107:{38,38}]
  wire  _GEN_767 = 7'h78 == reqIndex ? way1Age_120 : _GEN_766; // @[ICache.scala 107:{38,38}]
  wire  _GEN_768 = 7'h79 == reqIndex ? way1Age_121 : _GEN_767; // @[ICache.scala 107:{38,38}]
  wire  _GEN_769 = 7'h7a == reqIndex ? way1Age_122 : _GEN_768; // @[ICache.scala 107:{38,38}]
  wire  _GEN_770 = 7'h7b == reqIndex ? way1Age_123 : _GEN_769; // @[ICache.scala 107:{38,38}]
  wire  _GEN_771 = 7'h7c == reqIndex ? way1Age_124 : _GEN_770; // @[ICache.scala 107:{38,38}]
  wire  _GEN_772 = 7'h7d == reqIndex ? way1Age_125 : _GEN_771; // @[ICache.scala 107:{38,38}]
  wire  _GEN_773 = 7'h7e == reqIndex ? way1Age_126 : _GEN_772; // @[ICache.scala 107:{38,38}]
  wire  _GEN_774 = 7'h7f == reqIndex ? way1Age_127 : _GEN_773; // @[ICache.scala 107:{38,38}]
  wire  ageWay1En = ~_GEN_774 & sFillEn; // @[ICache.scala 107:47]
  wire  _GEN_2311 = 7'h0 == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1159 = 7'h0 == reqIndex | way0V_0; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2312 = 7'h1 == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1160 = 7'h1 == reqIndex | way0V_1; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2313 = 7'h2 == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1161 = 7'h2 == reqIndex | way0V_2; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2314 = 7'h3 == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1162 = 7'h3 == reqIndex | way0V_3; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2315 = 7'h4 == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1163 = 7'h4 == reqIndex | way0V_4; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2316 = 7'h5 == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1164 = 7'h5 == reqIndex | way0V_5; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2317 = 7'h6 == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1165 = 7'h6 == reqIndex | way0V_6; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2318 = 7'h7 == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1166 = 7'h7 == reqIndex | way0V_7; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2319 = 7'h8 == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1167 = 7'h8 == reqIndex | way0V_8; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2320 = 7'h9 == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1168 = 7'h9 == reqIndex | way0V_9; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2321 = 7'ha == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1169 = 7'ha == reqIndex | way0V_10; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2322 = 7'hb == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1170 = 7'hb == reqIndex | way0V_11; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2323 = 7'hc == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1171 = 7'hc == reqIndex | way0V_12; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2324 = 7'hd == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1172 = 7'hd == reqIndex | way0V_13; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2325 = 7'he == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1173 = 7'he == reqIndex | way0V_14; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2326 = 7'hf == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1174 = 7'hf == reqIndex | way0V_15; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2327 = 7'h10 == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1175 = 7'h10 == reqIndex | way0V_16; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2328 = 7'h11 == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1176 = 7'h11 == reqIndex | way0V_17; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2329 = 7'h12 == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1177 = 7'h12 == reqIndex | way0V_18; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2330 = 7'h13 == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1178 = 7'h13 == reqIndex | way0V_19; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2331 = 7'h14 == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1179 = 7'h14 == reqIndex | way0V_20; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2332 = 7'h15 == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1180 = 7'h15 == reqIndex | way0V_21; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2333 = 7'h16 == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1181 = 7'h16 == reqIndex | way0V_22; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2334 = 7'h17 == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1182 = 7'h17 == reqIndex | way0V_23; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2335 = 7'h18 == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1183 = 7'h18 == reqIndex | way0V_24; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2336 = 7'h19 == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1184 = 7'h19 == reqIndex | way0V_25; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2337 = 7'h1a == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1185 = 7'h1a == reqIndex | way0V_26; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2338 = 7'h1b == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1186 = 7'h1b == reqIndex | way0V_27; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2339 = 7'h1c == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1187 = 7'h1c == reqIndex | way0V_28; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2340 = 7'h1d == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1188 = 7'h1d == reqIndex | way0V_29; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2341 = 7'h1e == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1189 = 7'h1e == reqIndex | way0V_30; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2342 = 7'h1f == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1190 = 7'h1f == reqIndex | way0V_31; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2343 = 7'h20 == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1191 = 7'h20 == reqIndex | way0V_32; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2344 = 7'h21 == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1192 = 7'h21 == reqIndex | way0V_33; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2345 = 7'h22 == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1193 = 7'h22 == reqIndex | way0V_34; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2346 = 7'h23 == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1194 = 7'h23 == reqIndex | way0V_35; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2347 = 7'h24 == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1195 = 7'h24 == reqIndex | way0V_36; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2348 = 7'h25 == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1196 = 7'h25 == reqIndex | way0V_37; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2349 = 7'h26 == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1197 = 7'h26 == reqIndex | way0V_38; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2350 = 7'h27 == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1198 = 7'h27 == reqIndex | way0V_39; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2351 = 7'h28 == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1199 = 7'h28 == reqIndex | way0V_40; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2352 = 7'h29 == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1200 = 7'h29 == reqIndex | way0V_41; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2353 = 7'h2a == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1201 = 7'h2a == reqIndex | way0V_42; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2354 = 7'h2b == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1202 = 7'h2b == reqIndex | way0V_43; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2355 = 7'h2c == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1203 = 7'h2c == reqIndex | way0V_44; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2356 = 7'h2d == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1204 = 7'h2d == reqIndex | way0V_45; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2357 = 7'h2e == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1205 = 7'h2e == reqIndex | way0V_46; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2358 = 7'h2f == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1206 = 7'h2f == reqIndex | way0V_47; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2359 = 7'h30 == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1207 = 7'h30 == reqIndex | way0V_48; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2360 = 7'h31 == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1208 = 7'h31 == reqIndex | way0V_49; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2361 = 7'h32 == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1209 = 7'h32 == reqIndex | way0V_50; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2362 = 7'h33 == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1210 = 7'h33 == reqIndex | way0V_51; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2363 = 7'h34 == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1211 = 7'h34 == reqIndex | way0V_52; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2364 = 7'h35 == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1212 = 7'h35 == reqIndex | way0V_53; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2365 = 7'h36 == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1213 = 7'h36 == reqIndex | way0V_54; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2366 = 7'h37 == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1214 = 7'h37 == reqIndex | way0V_55; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2367 = 7'h38 == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1215 = 7'h38 == reqIndex | way0V_56; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2368 = 7'h39 == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1216 = 7'h39 == reqIndex | way0V_57; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2369 = 7'h3a == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1217 = 7'h3a == reqIndex | way0V_58; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2370 = 7'h3b == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1218 = 7'h3b == reqIndex | way0V_59; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2371 = 7'h3c == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1219 = 7'h3c == reqIndex | way0V_60; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2372 = 7'h3d == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1220 = 7'h3d == reqIndex | way0V_61; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2373 = 7'h3e == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1221 = 7'h3e == reqIndex | way0V_62; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2374 = 7'h3f == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1222 = 7'h3f == reqIndex | way0V_63; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2375 = 7'h40 == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1223 = 7'h40 == reqIndex | way0V_64; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2376 = 7'h41 == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1224 = 7'h41 == reqIndex | way0V_65; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2377 = 7'h42 == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1225 = 7'h42 == reqIndex | way0V_66; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2378 = 7'h43 == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1226 = 7'h43 == reqIndex | way0V_67; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2379 = 7'h44 == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1227 = 7'h44 == reqIndex | way0V_68; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2380 = 7'h45 == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1228 = 7'h45 == reqIndex | way0V_69; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2381 = 7'h46 == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1229 = 7'h46 == reqIndex | way0V_70; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2382 = 7'h47 == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1230 = 7'h47 == reqIndex | way0V_71; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2383 = 7'h48 == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1231 = 7'h48 == reqIndex | way0V_72; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2384 = 7'h49 == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1232 = 7'h49 == reqIndex | way0V_73; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2385 = 7'h4a == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1233 = 7'h4a == reqIndex | way0V_74; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2386 = 7'h4b == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1234 = 7'h4b == reqIndex | way0V_75; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2387 = 7'h4c == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1235 = 7'h4c == reqIndex | way0V_76; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2388 = 7'h4d == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1236 = 7'h4d == reqIndex | way0V_77; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2389 = 7'h4e == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1237 = 7'h4e == reqIndex | way0V_78; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2390 = 7'h4f == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1238 = 7'h4f == reqIndex | way0V_79; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2391 = 7'h50 == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1239 = 7'h50 == reqIndex | way0V_80; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2392 = 7'h51 == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1240 = 7'h51 == reqIndex | way0V_81; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2393 = 7'h52 == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1241 = 7'h52 == reqIndex | way0V_82; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2394 = 7'h53 == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1242 = 7'h53 == reqIndex | way0V_83; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2395 = 7'h54 == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1243 = 7'h54 == reqIndex | way0V_84; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2396 = 7'h55 == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1244 = 7'h55 == reqIndex | way0V_85; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2397 = 7'h56 == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1245 = 7'h56 == reqIndex | way0V_86; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2398 = 7'h57 == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1246 = 7'h57 == reqIndex | way0V_87; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2399 = 7'h58 == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1247 = 7'h58 == reqIndex | way0V_88; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2400 = 7'h59 == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1248 = 7'h59 == reqIndex | way0V_89; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2401 = 7'h5a == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1249 = 7'h5a == reqIndex | way0V_90; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2402 = 7'h5b == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1250 = 7'h5b == reqIndex | way0V_91; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2403 = 7'h5c == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1251 = 7'h5c == reqIndex | way0V_92; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2404 = 7'h5d == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1252 = 7'h5d == reqIndex | way0V_93; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2405 = 7'h5e == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1253 = 7'h5e == reqIndex | way0V_94; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2406 = 7'h5f == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1254 = 7'h5f == reqIndex | way0V_95; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2407 = 7'h60 == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1255 = 7'h60 == reqIndex | way0V_96; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2408 = 7'h61 == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1256 = 7'h61 == reqIndex | way0V_97; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2409 = 7'h62 == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1257 = 7'h62 == reqIndex | way0V_98; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2410 = 7'h63 == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1258 = 7'h63 == reqIndex | way0V_99; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2411 = 7'h64 == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1259 = 7'h64 == reqIndex | way0V_100; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2412 = 7'h65 == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1260 = 7'h65 == reqIndex | way0V_101; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2413 = 7'h66 == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1261 = 7'h66 == reqIndex | way0V_102; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2414 = 7'h67 == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1262 = 7'h67 == reqIndex | way0V_103; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2415 = 7'h68 == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1263 = 7'h68 == reqIndex | way0V_104; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2416 = 7'h69 == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1264 = 7'h69 == reqIndex | way0V_105; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2417 = 7'h6a == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1265 = 7'h6a == reqIndex | way0V_106; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2418 = 7'h6b == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1266 = 7'h6b == reqIndex | way0V_107; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2419 = 7'h6c == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1267 = 7'h6c == reqIndex | way0V_108; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2420 = 7'h6d == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1268 = 7'h6d == reqIndex | way0V_109; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2421 = 7'h6e == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1269 = 7'h6e == reqIndex | way0V_110; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2422 = 7'h6f == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1270 = 7'h6f == reqIndex | way0V_111; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2423 = 7'h70 == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1271 = 7'h70 == reqIndex | way0V_112; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2424 = 7'h71 == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1272 = 7'h71 == reqIndex | way0V_113; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2425 = 7'h72 == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1273 = 7'h72 == reqIndex | way0V_114; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2426 = 7'h73 == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1274 = 7'h73 == reqIndex | way0V_115; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2427 = 7'h74 == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1275 = 7'h74 == reqIndex | way0V_116; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2428 = 7'h75 == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1276 = 7'h75 == reqIndex | way0V_117; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2429 = 7'h76 == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1277 = 7'h76 == reqIndex | way0V_118; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2430 = 7'h77 == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1278 = 7'h77 == reqIndex | way0V_119; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2431 = 7'h78 == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1279 = 7'h78 == reqIndex | way0V_120; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2432 = 7'h79 == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1280 = 7'h79 == reqIndex | way0V_121; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2433 = 7'h7a == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1281 = 7'h7a == reqIndex | way0V_122; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2434 = 7'h7b == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1282 = 7'h7b == reqIndex | way0V_123; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2435 = 7'h7c == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1283 = 7'h7c == reqIndex | way0V_124; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2436 = 7'h7d == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1284 = 7'h7d == reqIndex | way0V_125; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2437 = 7'h7e == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1285 = 7'h7e == reqIndex | way0V_126; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_2438 = 7'h7f == reqIndex; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1286 = 7'h7f == reqIndex | way0V_127; // @[ICache.scala 116:{21,21} 27:22]
  wire  _GEN_1415 = _GEN_2311 | way1V_0; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1416 = _GEN_2312 | way1V_1; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1417 = _GEN_2313 | way1V_2; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1418 = _GEN_2314 | way1V_3; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1419 = _GEN_2315 | way1V_4; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1420 = _GEN_2316 | way1V_5; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1421 = _GEN_2317 | way1V_6; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1422 = _GEN_2318 | way1V_7; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1423 = _GEN_2319 | way1V_8; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1424 = _GEN_2320 | way1V_9; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1425 = _GEN_2321 | way1V_10; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1426 = _GEN_2322 | way1V_11; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1427 = _GEN_2323 | way1V_12; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1428 = _GEN_2324 | way1V_13; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1429 = _GEN_2325 | way1V_14; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1430 = _GEN_2326 | way1V_15; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1431 = _GEN_2327 | way1V_16; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1432 = _GEN_2328 | way1V_17; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1433 = _GEN_2329 | way1V_18; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1434 = _GEN_2330 | way1V_19; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1435 = _GEN_2331 | way1V_20; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1436 = _GEN_2332 | way1V_21; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1437 = _GEN_2333 | way1V_22; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1438 = _GEN_2334 | way1V_23; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1439 = _GEN_2335 | way1V_24; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1440 = _GEN_2336 | way1V_25; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1441 = _GEN_2337 | way1V_26; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1442 = _GEN_2338 | way1V_27; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1443 = _GEN_2339 | way1V_28; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1444 = _GEN_2340 | way1V_29; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1445 = _GEN_2341 | way1V_30; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1446 = _GEN_2342 | way1V_31; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1447 = _GEN_2343 | way1V_32; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1448 = _GEN_2344 | way1V_33; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1449 = _GEN_2345 | way1V_34; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1450 = _GEN_2346 | way1V_35; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1451 = _GEN_2347 | way1V_36; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1452 = _GEN_2348 | way1V_37; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1453 = _GEN_2349 | way1V_38; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1454 = _GEN_2350 | way1V_39; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1455 = _GEN_2351 | way1V_40; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1456 = _GEN_2352 | way1V_41; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1457 = _GEN_2353 | way1V_42; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1458 = _GEN_2354 | way1V_43; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1459 = _GEN_2355 | way1V_44; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1460 = _GEN_2356 | way1V_45; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1461 = _GEN_2357 | way1V_46; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1462 = _GEN_2358 | way1V_47; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1463 = _GEN_2359 | way1V_48; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1464 = _GEN_2360 | way1V_49; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1465 = _GEN_2361 | way1V_50; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1466 = _GEN_2362 | way1V_51; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1467 = _GEN_2363 | way1V_52; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1468 = _GEN_2364 | way1V_53; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1469 = _GEN_2365 | way1V_54; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1470 = _GEN_2366 | way1V_55; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1471 = _GEN_2367 | way1V_56; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1472 = _GEN_2368 | way1V_57; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1473 = _GEN_2369 | way1V_58; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1474 = _GEN_2370 | way1V_59; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1475 = _GEN_2371 | way1V_60; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1476 = _GEN_2372 | way1V_61; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1477 = _GEN_2373 | way1V_62; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1478 = _GEN_2374 | way1V_63; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1479 = _GEN_2375 | way1V_64; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1480 = _GEN_2376 | way1V_65; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1481 = _GEN_2377 | way1V_66; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1482 = _GEN_2378 | way1V_67; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1483 = _GEN_2379 | way1V_68; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1484 = _GEN_2380 | way1V_69; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1485 = _GEN_2381 | way1V_70; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1486 = _GEN_2382 | way1V_71; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1487 = _GEN_2383 | way1V_72; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1488 = _GEN_2384 | way1V_73; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1489 = _GEN_2385 | way1V_74; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1490 = _GEN_2386 | way1V_75; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1491 = _GEN_2387 | way1V_76; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1492 = _GEN_2388 | way1V_77; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1493 = _GEN_2389 | way1V_78; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1494 = _GEN_2390 | way1V_79; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1495 = _GEN_2391 | way1V_80; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1496 = _GEN_2392 | way1V_81; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1497 = _GEN_2393 | way1V_82; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1498 = _GEN_2394 | way1V_83; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1499 = _GEN_2395 | way1V_84; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1500 = _GEN_2396 | way1V_85; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1501 = _GEN_2397 | way1V_86; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1502 = _GEN_2398 | way1V_87; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1503 = _GEN_2399 | way1V_88; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1504 = _GEN_2400 | way1V_89; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1505 = _GEN_2401 | way1V_90; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1506 = _GEN_2402 | way1V_91; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1507 = _GEN_2403 | way1V_92; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1508 = _GEN_2404 | way1V_93; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1509 = _GEN_2405 | way1V_94; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1510 = _GEN_2406 | way1V_95; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1511 = _GEN_2407 | way1V_96; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1512 = _GEN_2408 | way1V_97; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1513 = _GEN_2409 | way1V_98; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1514 = _GEN_2410 | way1V_99; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1515 = _GEN_2411 | way1V_100; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1516 = _GEN_2412 | way1V_101; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1517 = _GEN_2413 | way1V_102; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1518 = _GEN_2414 | way1V_103; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1519 = _GEN_2415 | way1V_104; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1520 = _GEN_2416 | way1V_105; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1521 = _GEN_2417 | way1V_106; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1522 = _GEN_2418 | way1V_107; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1523 = _GEN_2419 | way1V_108; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1524 = _GEN_2420 | way1V_109; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1525 = _GEN_2421 | way1V_110; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1526 = _GEN_2422 | way1V_111; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1527 = _GEN_2423 | way1V_112; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1528 = _GEN_2424 | way1V_113; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1529 = _GEN_2425 | way1V_114; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1530 = _GEN_2426 | way1V_115; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1531 = _GEN_2427 | way1V_116; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1532 = _GEN_2428 | way1V_117; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1533 = _GEN_2429 | way1V_118; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1534 = _GEN_2430 | way1V_119; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1535 = _GEN_2431 | way1V_120; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1536 = _GEN_2432 | way1V_121; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1537 = _GEN_2433 | way1V_122; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1538 = _GEN_2434 | way1V_123; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1539 = _GEN_2435 | way1V_124; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1540 = _GEN_2436 | way1V_125; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1541 = _GEN_2437 | way1V_126; // @[ICache.scala 119:{21,21} 32:22]
  wire  _GEN_1542 = _GEN_2438 | way1V_127; // @[ICache.scala 119:{21,21} 32:22]
  S011HD1P_X32Y2D128 req ( // @[ICache.scala 51:19]
    .Q(req_Q),
    .CLK(req_CLK),
    .CEN(req_CEN),
    .WEN(req_WEN),
    .A(req_A),
    .D(req_D)
  );
  assign io_imem_inst_ready = sReadEn & cacheHitEn; // @[ICache.scala 88:28]
  assign io_imem_inst_read = 2'h3 == reqOff[3:2] ? rData[127:96] : _io_imem_inst_read_T_8; // @[Mux.scala 81:58]
  assign io_out_inst_valid = state == 2'h2; // @[ICache.scala 96:22]
  assign io_out_inst_addr = sAxiEn ? io_imem_inst_addr : 32'h0; // @[ICache.scala 99:23]
  assign req_CLK = clock; // @[ICache.scala 52:14]
  assign req_CEN = 1'h1; // @[ICache.scala 53:14]
  assign req_WEN = state == 2'h3; // @[ICache.scala 104:23]
  assign req_A = ~sFillEn ? cacheRIndex : cacheWIndex; // @[ICache.scala 55:20]
  assign req_D = cacheWData; // @[ICache.scala 56:14]
  always @(posedge clock) begin
    if (reset) begin // @[ICache.scala 22:27]
      cacheWData <= 128'h0; // @[ICache.scala 22:27]
    end else if (sAxiEn & io_out_inst_ready) begin // @[ICache.scala 101:20]
      cacheWData <= io_out_inst_read;
    end else begin
      cacheWData <= 128'h0;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_0 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_0 <= _GEN_1159;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_1 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_1 <= _GEN_1160;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_2 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_2 <= _GEN_1161;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_3 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_3 <= _GEN_1162;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_4 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_4 <= _GEN_1163;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_5 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_5 <= _GEN_1164;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_6 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_6 <= _GEN_1165;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_7 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_7 <= _GEN_1166;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_8 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_8 <= _GEN_1167;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_9 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_9 <= _GEN_1168;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_10 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_10 <= _GEN_1169;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_11 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_11 <= _GEN_1170;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_12 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_12 <= _GEN_1171;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_13 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_13 <= _GEN_1172;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_14 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_14 <= _GEN_1173;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_15 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_15 <= _GEN_1174;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_16 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_16 <= _GEN_1175;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_17 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_17 <= _GEN_1176;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_18 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_18 <= _GEN_1177;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_19 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_19 <= _GEN_1178;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_20 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_20 <= _GEN_1179;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_21 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_21 <= _GEN_1180;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_22 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_22 <= _GEN_1181;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_23 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_23 <= _GEN_1182;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_24 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_24 <= _GEN_1183;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_25 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_25 <= _GEN_1184;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_26 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_26 <= _GEN_1185;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_27 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_27 <= _GEN_1186;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_28 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_28 <= _GEN_1187;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_29 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_29 <= _GEN_1188;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_30 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_30 <= _GEN_1189;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_31 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_31 <= _GEN_1190;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_32 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_32 <= _GEN_1191;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_33 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_33 <= _GEN_1192;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_34 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_34 <= _GEN_1193;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_35 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_35 <= _GEN_1194;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_36 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_36 <= _GEN_1195;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_37 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_37 <= _GEN_1196;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_38 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_38 <= _GEN_1197;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_39 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_39 <= _GEN_1198;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_40 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_40 <= _GEN_1199;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_41 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_41 <= _GEN_1200;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_42 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_42 <= _GEN_1201;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_43 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_43 <= _GEN_1202;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_44 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_44 <= _GEN_1203;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_45 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_45 <= _GEN_1204;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_46 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_46 <= _GEN_1205;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_47 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_47 <= _GEN_1206;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_48 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_48 <= _GEN_1207;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_49 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_49 <= _GEN_1208;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_50 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_50 <= _GEN_1209;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_51 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_51 <= _GEN_1210;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_52 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_52 <= _GEN_1211;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_53 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_53 <= _GEN_1212;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_54 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_54 <= _GEN_1213;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_55 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_55 <= _GEN_1214;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_56 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_56 <= _GEN_1215;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_57 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_57 <= _GEN_1216;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_58 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_58 <= _GEN_1217;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_59 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_59 <= _GEN_1218;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_60 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_60 <= _GEN_1219;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_61 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_61 <= _GEN_1220;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_62 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_62 <= _GEN_1221;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_63 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_63 <= _GEN_1222;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_64 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_64 <= _GEN_1223;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_65 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_65 <= _GEN_1224;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_66 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_66 <= _GEN_1225;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_67 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_67 <= _GEN_1226;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_68 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_68 <= _GEN_1227;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_69 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_69 <= _GEN_1228;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_70 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_70 <= _GEN_1229;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_71 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_71 <= _GEN_1230;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_72 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_72 <= _GEN_1231;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_73 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_73 <= _GEN_1232;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_74 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_74 <= _GEN_1233;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_75 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_75 <= _GEN_1234;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_76 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_76 <= _GEN_1235;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_77 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_77 <= _GEN_1236;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_78 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_78 <= _GEN_1237;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_79 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_79 <= _GEN_1238;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_80 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_80 <= _GEN_1239;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_81 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_81 <= _GEN_1240;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_82 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_82 <= _GEN_1241;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_83 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_83 <= _GEN_1242;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_84 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_84 <= _GEN_1243;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_85 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_85 <= _GEN_1244;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_86 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_86 <= _GEN_1245;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_87 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_87 <= _GEN_1246;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_88 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_88 <= _GEN_1247;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_89 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_89 <= _GEN_1248;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_90 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_90 <= _GEN_1249;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_91 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_91 <= _GEN_1250;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_92 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_92 <= _GEN_1251;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_93 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_93 <= _GEN_1252;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_94 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_94 <= _GEN_1253;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_95 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_95 <= _GEN_1254;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_96 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_96 <= _GEN_1255;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_97 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_97 <= _GEN_1256;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_98 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_98 <= _GEN_1257;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_99 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_99 <= _GEN_1258;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_100 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_100 <= _GEN_1259;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_101 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_101 <= _GEN_1260;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_102 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_102 <= _GEN_1261;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_103 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_103 <= _GEN_1262;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_104 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_104 <= _GEN_1263;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_105 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_105 <= _GEN_1264;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_106 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_106 <= _GEN_1265;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_107 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_107 <= _GEN_1266;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_108 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_108 <= _GEN_1267;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_109 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_109 <= _GEN_1268;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_110 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_110 <= _GEN_1269;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_111 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_111 <= _GEN_1270;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_112 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_112 <= _GEN_1271;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_113 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_113 <= _GEN_1272;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_114 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_114 <= _GEN_1273;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_115 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_115 <= _GEN_1274;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_116 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_116 <= _GEN_1275;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_117 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_117 <= _GEN_1276;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_118 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_118 <= _GEN_1277;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_119 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_119 <= _GEN_1278;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_120 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_120 <= _GEN_1279;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_121 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_121 <= _GEN_1280;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_122 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_122 <= _GEN_1281;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_123 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_123 <= _GEN_1282;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_124 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_124 <= _GEN_1283;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_125 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_125 <= _GEN_1284;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_126 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_126 <= _GEN_1285;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_127 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      way0V_127 <= _GEN_1286;
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_0 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h0 == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_0 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_1 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h1 == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_1 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_2 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h2 == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_2 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_3 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h3 == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_3 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_4 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h4 == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_4 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_5 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h5 == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_5 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_6 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h6 == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_6 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_7 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h7 == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_7 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_8 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h8 == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_8 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_9 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h9 == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_9 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_10 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'ha == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_10 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_11 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'hb == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_11 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_12 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'hc == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_12 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_13 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'hd == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_13 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_14 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'he == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_14 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_15 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'hf == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_15 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_16 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h10 == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_16 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_17 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h11 == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_17 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_18 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h12 == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_18 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_19 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h13 == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_19 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_20 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h14 == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_20 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_21 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h15 == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_21 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_22 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h16 == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_22 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_23 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h17 == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_23 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_24 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h18 == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_24 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_25 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h19 == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_25 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_26 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h1a == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_26 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_27 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h1b == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_27 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_28 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h1c == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_28 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_29 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h1d == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_29 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_30 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h1e == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_30 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_31 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h1f == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_31 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_32 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h20 == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_32 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_33 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h21 == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_33 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_34 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h22 == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_34 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_35 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h23 == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_35 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_36 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h24 == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_36 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_37 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h25 == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_37 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_38 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h26 == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_38 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_39 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h27 == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_39 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_40 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h28 == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_40 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_41 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h29 == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_41 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_42 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h2a == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_42 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_43 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h2b == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_43 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_44 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h2c == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_44 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_45 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h2d == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_45 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_46 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h2e == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_46 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_47 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h2f == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_47 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_48 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h30 == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_48 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_49 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h31 == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_49 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_50 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h32 == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_50 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_51 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h33 == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_51 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_52 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h34 == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_52 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_53 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h35 == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_53 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_54 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h36 == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_54 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_55 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h37 == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_55 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_56 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h38 == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_56 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_57 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h39 == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_57 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_58 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h3a == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_58 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_59 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h3b == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_59 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_60 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h3c == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_60 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_61 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h3d == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_61 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_62 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h3e == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_62 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_63 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h3f == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_63 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_64 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h40 == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_64 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_65 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h41 == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_65 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_66 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h42 == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_66 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_67 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h43 == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_67 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_68 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h44 == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_68 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_69 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h45 == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_69 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_70 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h46 == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_70 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_71 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h47 == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_71 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_72 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h48 == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_72 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_73 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h49 == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_73 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_74 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h4a == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_74 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_75 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h4b == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_75 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_76 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h4c == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_76 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_77 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h4d == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_77 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_78 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h4e == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_78 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_79 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h4f == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_79 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_80 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h50 == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_80 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_81 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h51 == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_81 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_82 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h52 == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_82 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_83 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h53 == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_83 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_84 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h54 == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_84 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_85 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h55 == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_85 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_86 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h56 == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_86 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_87 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h57 == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_87 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_88 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h58 == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_88 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_89 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h59 == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_89 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_90 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h5a == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_90 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_91 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h5b == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_91 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_92 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h5c == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_92 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_93 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h5d == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_93 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_94 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h5e == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_94 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_95 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h5f == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_95 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_96 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h60 == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_96 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_97 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h61 == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_97 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_98 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h62 == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_98 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_99 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h63 == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_99 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_100 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h64 == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_100 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_101 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h65 == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_101 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_102 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h66 == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_102 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_103 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h67 == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_103 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_104 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h68 == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_104 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_105 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h69 == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_105 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_106 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h6a == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_106 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_107 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h6b == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_107 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_108 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h6c == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_108 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_109 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h6d == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_109 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_110 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h6e == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_110 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_111 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h6f == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_111 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_112 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h70 == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_112 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_113 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h71 == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_113 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_114 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h72 == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_114 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_115 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h73 == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_115 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_116 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h74 == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_116 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_117 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h75 == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_117 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_118 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h76 == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_118 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_119 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h77 == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_119 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_120 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h78 == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_120 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_121 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h79 == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_121 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_122 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h7a == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_122 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_123 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h7b == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_123 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_124 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h7c == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_124 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_125 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h7d == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_125 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_126 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h7e == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_126 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_127 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 114:19]
      if (7'h7f == reqIndex) begin // @[ICache.scala 115:23]
        way0Tag_127 <= reqTag; // @[ICache.scala 115:23]
      end
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_0 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h0 == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_0 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_1 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h1 == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_1 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_2 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h2 == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_2 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_3 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h3 == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_3 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_4 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h4 == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_4 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_5 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h5 == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_5 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_6 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h6 == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_6 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_7 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h7 == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_7 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_8 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h8 == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_8 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_9 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h9 == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_9 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_10 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'ha == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_10 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_11 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'hb == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_11 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_12 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'hc == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_12 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_13 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'hd == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_13 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_14 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'he == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_14 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_15 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'hf == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_15 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_16 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h10 == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_16 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_17 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h11 == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_17 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_18 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h12 == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_18 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_19 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h13 == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_19 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_20 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h14 == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_20 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_21 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h15 == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_21 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_22 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h16 == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_22 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_23 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h17 == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_23 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_24 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h18 == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_24 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_25 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h19 == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_25 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_26 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h1a == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_26 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_27 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h1b == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_27 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_28 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h1c == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_28 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_29 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h1d == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_29 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_30 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h1e == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_30 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_31 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h1f == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_31 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_32 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h20 == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_32 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_33 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h21 == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_33 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_34 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h22 == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_34 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_35 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h23 == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_35 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_36 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h24 == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_36 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_37 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h25 == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_37 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_38 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h26 == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_38 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_39 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h27 == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_39 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_40 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h28 == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_40 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_41 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h29 == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_41 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_42 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h2a == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_42 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_43 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h2b == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_43 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_44 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h2c == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_44 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_45 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h2d == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_45 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_46 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h2e == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_46 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_47 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h2f == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_47 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_48 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h30 == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_48 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_49 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h31 == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_49 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_50 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h32 == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_50 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_51 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h33 == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_51 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_52 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h34 == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_52 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_53 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h35 == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_53 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_54 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h36 == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_54 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_55 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h37 == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_55 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_56 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h38 == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_56 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_57 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h39 == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_57 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_58 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h3a == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_58 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_59 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h3b == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_59 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_60 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h3c == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_60 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_61 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h3d == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_61 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_62 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h3e == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_62 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_63 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h3f == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_63 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_64 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h40 == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_64 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_65 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h41 == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_65 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_66 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h42 == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_66 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_67 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h43 == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_67 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_68 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h44 == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_68 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_69 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h45 == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_69 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_70 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h46 == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_70 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_71 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h47 == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_71 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_72 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h48 == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_72 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_73 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h49 == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_73 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_74 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h4a == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_74 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_75 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h4b == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_75 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_76 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h4c == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_76 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_77 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h4d == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_77 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_78 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h4e == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_78 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_79 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h4f == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_79 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_80 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h50 == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_80 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_81 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h51 == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_81 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_82 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h52 == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_82 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_83 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h53 == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_83 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_84 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h54 == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_84 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_85 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h55 == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_85 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_86 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h56 == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_86 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_87 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h57 == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_87 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_88 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h58 == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_88 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_89 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h59 == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_89 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_90 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h5a == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_90 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_91 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h5b == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_91 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_92 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h5c == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_92 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_93 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h5d == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_93 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_94 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h5e == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_94 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_95 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h5f == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_95 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_96 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h60 == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_96 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_97 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h61 == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_97 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_98 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h62 == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_98 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_99 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h63 == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_99 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_100 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h64 == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_100 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_101 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h65 == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_101 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_102 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h66 == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_102 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_103 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h67 == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_103 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_104 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h68 == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_104 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_105 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h69 == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_105 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_106 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h6a == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_106 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_107 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h6b == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_107 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_108 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h6c == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_108 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_109 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h6d == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_109 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_110 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h6e == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_110 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_111 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h6f == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_111 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_112 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h70 == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_112 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_113 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h71 == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_113 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_114 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h72 == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_114 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_115 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h73 == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_115 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_116 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h74 == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_116 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_117 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h75 == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_117 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_118 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h76 == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_118 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_119 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h77 == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_119 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_120 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h78 == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_120 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_121 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h79 == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_121 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_122 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h7a == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_122 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_123 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h7b == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_123 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_124 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h7c == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_124 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_125 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h7d == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_125 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_126 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h7e == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_126 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_127 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h7f == reqIndex) begin // @[ICache.scala 109:21]
      way0Age_127 <= ageWay0En; // @[ICache.scala 109:21]
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_0 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_0 <= _GEN_1415;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_1 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_1 <= _GEN_1416;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_2 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_2 <= _GEN_1417;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_3 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_3 <= _GEN_1418;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_4 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_4 <= _GEN_1419;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_5 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_5 <= _GEN_1420;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_6 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_6 <= _GEN_1421;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_7 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_7 <= _GEN_1422;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_8 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_8 <= _GEN_1423;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_9 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_9 <= _GEN_1424;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_10 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_10 <= _GEN_1425;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_11 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_11 <= _GEN_1426;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_12 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_12 <= _GEN_1427;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_13 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_13 <= _GEN_1428;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_14 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_14 <= _GEN_1429;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_15 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_15 <= _GEN_1430;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_16 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_16 <= _GEN_1431;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_17 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_17 <= _GEN_1432;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_18 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_18 <= _GEN_1433;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_19 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_19 <= _GEN_1434;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_20 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_20 <= _GEN_1435;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_21 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_21 <= _GEN_1436;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_22 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_22 <= _GEN_1437;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_23 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_23 <= _GEN_1438;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_24 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_24 <= _GEN_1439;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_25 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_25 <= _GEN_1440;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_26 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_26 <= _GEN_1441;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_27 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_27 <= _GEN_1442;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_28 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_28 <= _GEN_1443;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_29 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_29 <= _GEN_1444;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_30 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_30 <= _GEN_1445;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_31 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_31 <= _GEN_1446;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_32 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_32 <= _GEN_1447;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_33 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_33 <= _GEN_1448;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_34 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_34 <= _GEN_1449;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_35 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_35 <= _GEN_1450;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_36 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_36 <= _GEN_1451;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_37 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_37 <= _GEN_1452;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_38 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_38 <= _GEN_1453;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_39 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_39 <= _GEN_1454;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_40 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_40 <= _GEN_1455;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_41 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_41 <= _GEN_1456;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_42 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_42 <= _GEN_1457;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_43 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_43 <= _GEN_1458;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_44 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_44 <= _GEN_1459;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_45 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_45 <= _GEN_1460;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_46 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_46 <= _GEN_1461;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_47 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_47 <= _GEN_1462;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_48 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_48 <= _GEN_1463;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_49 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_49 <= _GEN_1464;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_50 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_50 <= _GEN_1465;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_51 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_51 <= _GEN_1466;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_52 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_52 <= _GEN_1467;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_53 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_53 <= _GEN_1468;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_54 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_54 <= _GEN_1469;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_55 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_55 <= _GEN_1470;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_56 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_56 <= _GEN_1471;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_57 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_57 <= _GEN_1472;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_58 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_58 <= _GEN_1473;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_59 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_59 <= _GEN_1474;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_60 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_60 <= _GEN_1475;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_61 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_61 <= _GEN_1476;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_62 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_62 <= _GEN_1477;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_63 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_63 <= _GEN_1478;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_64 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_64 <= _GEN_1479;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_65 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_65 <= _GEN_1480;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_66 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_66 <= _GEN_1481;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_67 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_67 <= _GEN_1482;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_68 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_68 <= _GEN_1483;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_69 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_69 <= _GEN_1484;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_70 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_70 <= _GEN_1485;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_71 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_71 <= _GEN_1486;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_72 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_72 <= _GEN_1487;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_73 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_73 <= _GEN_1488;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_74 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_74 <= _GEN_1489;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_75 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_75 <= _GEN_1490;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_76 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_76 <= _GEN_1491;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_77 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_77 <= _GEN_1492;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_78 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_78 <= _GEN_1493;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_79 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_79 <= _GEN_1494;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_80 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_80 <= _GEN_1495;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_81 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_81 <= _GEN_1496;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_82 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_82 <= _GEN_1497;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_83 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_83 <= _GEN_1498;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_84 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_84 <= _GEN_1499;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_85 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_85 <= _GEN_1500;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_86 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_86 <= _GEN_1501;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_87 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_87 <= _GEN_1502;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_88 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_88 <= _GEN_1503;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_89 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_89 <= _GEN_1504;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_90 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_90 <= _GEN_1505;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_91 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_91 <= _GEN_1506;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_92 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_92 <= _GEN_1507;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_93 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_93 <= _GEN_1508;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_94 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_94 <= _GEN_1509;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_95 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_95 <= _GEN_1510;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_96 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_96 <= _GEN_1511;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_97 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_97 <= _GEN_1512;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_98 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_98 <= _GEN_1513;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_99 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_99 <= _GEN_1514;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_100 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_100 <= _GEN_1515;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_101 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_101 <= _GEN_1516;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_102 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_102 <= _GEN_1517;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_103 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_103 <= _GEN_1518;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_104 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_104 <= _GEN_1519;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_105 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_105 <= _GEN_1520;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_106 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_106 <= _GEN_1521;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_107 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_107 <= _GEN_1522;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_108 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_108 <= _GEN_1523;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_109 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_109 <= _GEN_1524;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_110 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_110 <= _GEN_1525;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_111 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_111 <= _GEN_1526;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_112 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_112 <= _GEN_1527;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_113 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_113 <= _GEN_1528;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_114 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_114 <= _GEN_1529;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_115 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_115 <= _GEN_1530;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_116 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_116 <= _GEN_1531;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_117 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_117 <= _GEN_1532;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_118 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_118 <= _GEN_1533;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_119 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_119 <= _GEN_1534;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_120 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_120 <= _GEN_1535;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_121 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_121 <= _GEN_1536;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_122 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_122 <= _GEN_1537;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_123 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_123 <= _GEN_1538;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_124 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_124 <= _GEN_1539;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_125 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_125 <= _GEN_1540;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_126 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_126 <= _GEN_1541;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_127 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        way1V_127 <= _GEN_1542;
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_0 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h0 == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_0 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_1 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h1 == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_1 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_2 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h2 == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_2 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_3 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h3 == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_3 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_4 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h4 == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_4 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_5 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h5 == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_5 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_6 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h6 == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_6 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_7 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h7 == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_7 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_8 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h8 == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_8 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_9 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h9 == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_9 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_10 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'ha == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_10 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_11 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'hb == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_11 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_12 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'hc == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_12 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_13 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'hd == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_13 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_14 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'he == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_14 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_15 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'hf == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_15 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_16 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h10 == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_16 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_17 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h11 == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_17 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_18 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h12 == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_18 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_19 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h13 == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_19 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_20 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h14 == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_20 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_21 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h15 == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_21 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_22 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h16 == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_22 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_23 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h17 == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_23 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_24 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h18 == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_24 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_25 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h19 == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_25 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_26 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h1a == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_26 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_27 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h1b == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_27 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_28 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h1c == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_28 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_29 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h1d == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_29 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_30 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h1e == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_30 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_31 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h1f == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_31 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_32 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h20 == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_32 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_33 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h21 == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_33 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_34 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h22 == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_34 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_35 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h23 == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_35 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_36 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h24 == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_36 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_37 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h25 == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_37 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_38 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h26 == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_38 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_39 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h27 == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_39 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_40 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h28 == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_40 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_41 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h29 == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_41 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_42 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h2a == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_42 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_43 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h2b == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_43 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_44 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h2c == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_44 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_45 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h2d == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_45 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_46 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h2e == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_46 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_47 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h2f == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_47 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_48 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h30 == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_48 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_49 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h31 == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_49 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_50 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h32 == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_50 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_51 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h33 == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_51 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_52 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h34 == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_52 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_53 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h35 == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_53 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_54 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h36 == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_54 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_55 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h37 == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_55 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_56 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h38 == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_56 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_57 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h39 == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_57 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_58 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h3a == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_58 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_59 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h3b == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_59 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_60 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h3c == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_60 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_61 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h3d == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_61 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_62 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h3e == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_62 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_63 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h3f == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_63 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_64 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h40 == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_64 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_65 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h41 == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_65 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_66 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h42 == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_66 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_67 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h43 == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_67 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_68 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h44 == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_68 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_69 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h45 == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_69 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_70 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h46 == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_70 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_71 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h47 == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_71 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_72 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h48 == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_72 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_73 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h49 == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_73 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_74 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h4a == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_74 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_75 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h4b == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_75 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_76 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h4c == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_76 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_77 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h4d == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_77 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_78 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h4e == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_78 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_79 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h4f == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_79 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_80 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h50 == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_80 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_81 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h51 == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_81 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_82 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h52 == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_82 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_83 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h53 == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_83 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_84 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h54 == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_84 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_85 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h55 == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_85 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_86 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h56 == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_86 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_87 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h57 == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_87 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_88 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h58 == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_88 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_89 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h59 == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_89 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_90 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h5a == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_90 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_91 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h5b == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_91 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_92 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h5c == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_92 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_93 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h5d == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_93 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_94 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h5e == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_94 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_95 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h5f == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_95 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_96 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h60 == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_96 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_97 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h61 == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_97 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_98 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h62 == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_98 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_99 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h63 == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_99 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_100 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h64 == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_100 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_101 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h65 == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_101 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_102 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h66 == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_102 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_103 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h67 == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_103 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_104 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h68 == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_104 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_105 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h69 == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_105 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_106 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h6a == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_106 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_107 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h6b == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_107 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_108 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h6c == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_108 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_109 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h6d == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_109 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_110 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h6e == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_110 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_111 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h6f == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_111 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_112 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h70 == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_112 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_113 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h71 == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_113 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_114 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h72 == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_114 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_115 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h73 == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_115 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_116 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h74 == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_116 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_117 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h75 == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_117 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_118 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h76 == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_118 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_119 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h77 == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_119 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_120 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h78 == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_120 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_121 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h79 == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_121 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_122 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h7a == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_122 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_123 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h7b == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_123 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_124 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h7c == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_124 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_125 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h7d == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_125 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_126 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h7e == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_126 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_127 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 114:19]
      if (ageWay1En) begin // @[ICache.scala 117:26]
        if (7'h7f == reqIndex) begin // @[ICache.scala 118:23]
          way1Tag_127 <= reqTag; // @[ICache.scala 118:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_0 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h0 == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_0 <= 1'h0;
      end else begin
        way1Age_0 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_1 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h1 == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_1 <= 1'h0;
      end else begin
        way1Age_1 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_2 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h2 == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_2 <= 1'h0;
      end else begin
        way1Age_2 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_3 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h3 == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_3 <= 1'h0;
      end else begin
        way1Age_3 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_4 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h4 == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_4 <= 1'h0;
      end else begin
        way1Age_4 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_5 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h5 == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_5 <= 1'h0;
      end else begin
        way1Age_5 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_6 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h6 == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_6 <= 1'h0;
      end else begin
        way1Age_6 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_7 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h7 == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_7 <= 1'h0;
      end else begin
        way1Age_7 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_8 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h8 == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_8 <= 1'h0;
      end else begin
        way1Age_8 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_9 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h9 == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_9 <= 1'h0;
      end else begin
        way1Age_9 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_10 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'ha == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_10 <= 1'h0;
      end else begin
        way1Age_10 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_11 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'hb == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_11 <= 1'h0;
      end else begin
        way1Age_11 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_12 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'hc == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_12 <= 1'h0;
      end else begin
        way1Age_12 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_13 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'hd == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_13 <= 1'h0;
      end else begin
        way1Age_13 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_14 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'he == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_14 <= 1'h0;
      end else begin
        way1Age_14 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_15 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'hf == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_15 <= 1'h0;
      end else begin
        way1Age_15 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_16 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h10 == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_16 <= 1'h0;
      end else begin
        way1Age_16 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_17 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h11 == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_17 <= 1'h0;
      end else begin
        way1Age_17 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_18 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h12 == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_18 <= 1'h0;
      end else begin
        way1Age_18 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_19 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h13 == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_19 <= 1'h0;
      end else begin
        way1Age_19 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_20 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h14 == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_20 <= 1'h0;
      end else begin
        way1Age_20 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_21 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h15 == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_21 <= 1'h0;
      end else begin
        way1Age_21 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_22 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h16 == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_22 <= 1'h0;
      end else begin
        way1Age_22 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_23 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h17 == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_23 <= 1'h0;
      end else begin
        way1Age_23 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_24 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h18 == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_24 <= 1'h0;
      end else begin
        way1Age_24 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_25 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h19 == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_25 <= 1'h0;
      end else begin
        way1Age_25 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_26 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h1a == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_26 <= 1'h0;
      end else begin
        way1Age_26 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_27 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h1b == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_27 <= 1'h0;
      end else begin
        way1Age_27 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_28 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h1c == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_28 <= 1'h0;
      end else begin
        way1Age_28 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_29 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h1d == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_29 <= 1'h0;
      end else begin
        way1Age_29 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_30 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h1e == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_30 <= 1'h0;
      end else begin
        way1Age_30 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_31 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h1f == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_31 <= 1'h0;
      end else begin
        way1Age_31 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_32 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h20 == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_32 <= 1'h0;
      end else begin
        way1Age_32 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_33 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h21 == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_33 <= 1'h0;
      end else begin
        way1Age_33 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_34 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h22 == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_34 <= 1'h0;
      end else begin
        way1Age_34 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_35 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h23 == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_35 <= 1'h0;
      end else begin
        way1Age_35 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_36 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h24 == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_36 <= 1'h0;
      end else begin
        way1Age_36 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_37 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h25 == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_37 <= 1'h0;
      end else begin
        way1Age_37 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_38 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h26 == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_38 <= 1'h0;
      end else begin
        way1Age_38 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_39 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h27 == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_39 <= 1'h0;
      end else begin
        way1Age_39 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_40 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h28 == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_40 <= 1'h0;
      end else begin
        way1Age_40 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_41 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h29 == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_41 <= 1'h0;
      end else begin
        way1Age_41 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_42 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h2a == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_42 <= 1'h0;
      end else begin
        way1Age_42 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_43 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h2b == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_43 <= 1'h0;
      end else begin
        way1Age_43 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_44 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h2c == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_44 <= 1'h0;
      end else begin
        way1Age_44 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_45 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h2d == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_45 <= 1'h0;
      end else begin
        way1Age_45 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_46 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h2e == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_46 <= 1'h0;
      end else begin
        way1Age_46 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_47 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h2f == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_47 <= 1'h0;
      end else begin
        way1Age_47 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_48 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h30 == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_48 <= 1'h0;
      end else begin
        way1Age_48 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_49 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h31 == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_49 <= 1'h0;
      end else begin
        way1Age_49 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_50 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h32 == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_50 <= 1'h0;
      end else begin
        way1Age_50 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_51 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h33 == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_51 <= 1'h0;
      end else begin
        way1Age_51 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_52 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h34 == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_52 <= 1'h0;
      end else begin
        way1Age_52 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_53 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h35 == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_53 <= 1'h0;
      end else begin
        way1Age_53 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_54 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h36 == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_54 <= 1'h0;
      end else begin
        way1Age_54 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_55 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h37 == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_55 <= 1'h0;
      end else begin
        way1Age_55 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_56 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h38 == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_56 <= 1'h0;
      end else begin
        way1Age_56 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_57 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h39 == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_57 <= 1'h0;
      end else begin
        way1Age_57 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_58 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h3a == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_58 <= 1'h0;
      end else begin
        way1Age_58 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_59 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h3b == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_59 <= 1'h0;
      end else begin
        way1Age_59 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_60 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h3c == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_60 <= 1'h0;
      end else begin
        way1Age_60 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_61 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h3d == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_61 <= 1'h0;
      end else begin
        way1Age_61 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_62 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h3e == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_62 <= 1'h0;
      end else begin
        way1Age_62 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_63 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h3f == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_63 <= 1'h0;
      end else begin
        way1Age_63 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_64 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h40 == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_64 <= 1'h0;
      end else begin
        way1Age_64 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_65 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h41 == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_65 <= 1'h0;
      end else begin
        way1Age_65 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_66 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h42 == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_66 <= 1'h0;
      end else begin
        way1Age_66 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_67 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h43 == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_67 <= 1'h0;
      end else begin
        way1Age_67 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_68 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h44 == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_68 <= 1'h0;
      end else begin
        way1Age_68 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_69 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h45 == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_69 <= 1'h0;
      end else begin
        way1Age_69 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_70 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h46 == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_70 <= 1'h0;
      end else begin
        way1Age_70 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_71 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h47 == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_71 <= 1'h0;
      end else begin
        way1Age_71 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_72 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h48 == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_72 <= 1'h0;
      end else begin
        way1Age_72 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_73 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h49 == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_73 <= 1'h0;
      end else begin
        way1Age_73 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_74 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h4a == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_74 <= 1'h0;
      end else begin
        way1Age_74 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_75 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h4b == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_75 <= 1'h0;
      end else begin
        way1Age_75 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_76 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h4c == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_76 <= 1'h0;
      end else begin
        way1Age_76 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_77 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h4d == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_77 <= 1'h0;
      end else begin
        way1Age_77 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_78 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h4e == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_78 <= 1'h0;
      end else begin
        way1Age_78 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_79 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h4f == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_79 <= 1'h0;
      end else begin
        way1Age_79 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_80 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h50 == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_80 <= 1'h0;
      end else begin
        way1Age_80 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_81 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h51 == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_81 <= 1'h0;
      end else begin
        way1Age_81 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_82 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h52 == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_82 <= 1'h0;
      end else begin
        way1Age_82 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_83 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h53 == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_83 <= 1'h0;
      end else begin
        way1Age_83 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_84 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h54 == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_84 <= 1'h0;
      end else begin
        way1Age_84 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_85 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h55 == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_85 <= 1'h0;
      end else begin
        way1Age_85 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_86 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h56 == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_86 <= 1'h0;
      end else begin
        way1Age_86 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_87 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h57 == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_87 <= 1'h0;
      end else begin
        way1Age_87 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_88 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h58 == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_88 <= 1'h0;
      end else begin
        way1Age_88 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_89 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h59 == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_89 <= 1'h0;
      end else begin
        way1Age_89 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_90 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h5a == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_90 <= 1'h0;
      end else begin
        way1Age_90 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_91 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h5b == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_91 <= 1'h0;
      end else begin
        way1Age_91 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_92 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h5c == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_92 <= 1'h0;
      end else begin
        way1Age_92 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_93 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h5d == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_93 <= 1'h0;
      end else begin
        way1Age_93 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_94 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h5e == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_94 <= 1'h0;
      end else begin
        way1Age_94 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_95 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h5f == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_95 <= 1'h0;
      end else begin
        way1Age_95 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_96 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h60 == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_96 <= 1'h0;
      end else begin
        way1Age_96 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_97 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h61 == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_97 <= 1'h0;
      end else begin
        way1Age_97 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_98 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h62 == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_98 <= 1'h0;
      end else begin
        way1Age_98 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_99 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h63 == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_99 <= 1'h0;
      end else begin
        way1Age_99 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_100 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h64 == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_100 <= 1'h0;
      end else begin
        way1Age_100 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_101 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h65 == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_101 <= 1'h0;
      end else begin
        way1Age_101 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_102 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h66 == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_102 <= 1'h0;
      end else begin
        way1Age_102 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_103 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h67 == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_103 <= 1'h0;
      end else begin
        way1Age_103 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_104 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h68 == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_104 <= 1'h0;
      end else begin
        way1Age_104 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_105 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h69 == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_105 <= 1'h0;
      end else begin
        way1Age_105 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_106 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h6a == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_106 <= 1'h0;
      end else begin
        way1Age_106 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_107 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h6b == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_107 <= 1'h0;
      end else begin
        way1Age_107 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_108 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h6c == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_108 <= 1'h0;
      end else begin
        way1Age_108 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_109 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h6d == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_109 <= 1'h0;
      end else begin
        way1Age_109 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_110 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h6e == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_110 <= 1'h0;
      end else begin
        way1Age_110 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_111 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h6f == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_111 <= 1'h0;
      end else begin
        way1Age_111 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_112 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h70 == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_112 <= 1'h0;
      end else begin
        way1Age_112 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_113 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h71 == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_113 <= 1'h0;
      end else begin
        way1Age_113 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_114 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h72 == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_114 <= 1'h0;
      end else begin
        way1Age_114 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_115 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h73 == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_115 <= 1'h0;
      end else begin
        way1Age_115 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_116 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h74 == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_116 <= 1'h0;
      end else begin
        way1Age_116 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_117 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h75 == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_117 <= 1'h0;
      end else begin
        way1Age_117 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_118 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h76 == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_118 <= 1'h0;
      end else begin
        way1Age_118 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_119 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h77 == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_119 <= 1'h0;
      end else begin
        way1Age_119 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_120 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h78 == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_120 <= 1'h0;
      end else begin
        way1Age_120 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_121 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h79 == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_121 <= 1'h0;
      end else begin
        way1Age_121 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_122 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h7a == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_122 <= 1'h0;
      end else begin
        way1Age_122 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_123 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h7b == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_123 <= 1'h0;
      end else begin
        way1Age_123 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_124 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h7c == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_124 <= 1'h0;
      end else begin
        way1Age_124 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_125 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h7d == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_125 <= 1'h0;
      end else begin
        way1Age_125 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_126 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h7e == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_126 <= 1'h0;
      end else begin
        way1Age_126 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_127 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h7f == reqIndex) begin // @[ICache.scala 110:21]
      if (ageWay0En) begin // @[ICache.scala 108:25]
        way1Age_127 <= 1'h0;
      end else begin
        way1Age_127 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 38:22]
      state <= 2'h0; // @[ICache.scala 38:22]
    end else if (2'h0 == state) begin // @[ICache.scala 60:17]
      if (io_imem_inst_valid) begin // @[ICache.scala 62:27]
        state <= 2'h1; // @[ICache.scala 63:15]
      end
    end else if (2'h1 == state) begin // @[ICache.scala 60:17]
      if (cacheHitEn) begin // @[ICache.scala 68:24]
        state <= 2'h0; // @[ICache.scala 69:15]
      end else begin
        state <= 2'h2; // @[ICache.scala 71:15]
      end
    end else if (2'h2 == state) begin // @[ICache.scala 60:17]
      state <= _GEN_514;
    end else begin
      state <= _GEN_515;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {4{`RANDOM}};
  cacheWData = _RAND_0[127:0];
  _RAND_1 = {1{`RANDOM}};
  way0V_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  way0V_1 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  way0V_2 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  way0V_3 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  way0V_4 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  way0V_5 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  way0V_6 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  way0V_7 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  way0V_8 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  way0V_9 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  way0V_10 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  way0V_11 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  way0V_12 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  way0V_13 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  way0V_14 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  way0V_15 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  way0V_16 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  way0V_17 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  way0V_18 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  way0V_19 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  way0V_20 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  way0V_21 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  way0V_22 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  way0V_23 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  way0V_24 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  way0V_25 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  way0V_26 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  way0V_27 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  way0V_28 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  way0V_29 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  way0V_30 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  way0V_31 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  way0V_32 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  way0V_33 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  way0V_34 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  way0V_35 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  way0V_36 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  way0V_37 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  way0V_38 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  way0V_39 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  way0V_40 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  way0V_41 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  way0V_42 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  way0V_43 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  way0V_44 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  way0V_45 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  way0V_46 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  way0V_47 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  way0V_48 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  way0V_49 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  way0V_50 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  way0V_51 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  way0V_52 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  way0V_53 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  way0V_54 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  way0V_55 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  way0V_56 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  way0V_57 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  way0V_58 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  way0V_59 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  way0V_60 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  way0V_61 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  way0V_62 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  way0V_63 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  way0V_64 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  way0V_65 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  way0V_66 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  way0V_67 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  way0V_68 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  way0V_69 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  way0V_70 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  way0V_71 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  way0V_72 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  way0V_73 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  way0V_74 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  way0V_75 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  way0V_76 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  way0V_77 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  way0V_78 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  way0V_79 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  way0V_80 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  way0V_81 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  way0V_82 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  way0V_83 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  way0V_84 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  way0V_85 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  way0V_86 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  way0V_87 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  way0V_88 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  way0V_89 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  way0V_90 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  way0V_91 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  way0V_92 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  way0V_93 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  way0V_94 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  way0V_95 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  way0V_96 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  way0V_97 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  way0V_98 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  way0V_99 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  way0V_100 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  way0V_101 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  way0V_102 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  way0V_103 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  way0V_104 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  way0V_105 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  way0V_106 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  way0V_107 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  way0V_108 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  way0V_109 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  way0V_110 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  way0V_111 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  way0V_112 = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  way0V_113 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  way0V_114 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  way0V_115 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  way0V_116 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  way0V_117 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  way0V_118 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  way0V_119 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  way0V_120 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  way0V_121 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  way0V_122 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  way0V_123 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  way0V_124 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  way0V_125 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  way0V_126 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  way0V_127 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  way0Tag_0 = _RAND_129[20:0];
  _RAND_130 = {1{`RANDOM}};
  way0Tag_1 = _RAND_130[20:0];
  _RAND_131 = {1{`RANDOM}};
  way0Tag_2 = _RAND_131[20:0];
  _RAND_132 = {1{`RANDOM}};
  way0Tag_3 = _RAND_132[20:0];
  _RAND_133 = {1{`RANDOM}};
  way0Tag_4 = _RAND_133[20:0];
  _RAND_134 = {1{`RANDOM}};
  way0Tag_5 = _RAND_134[20:0];
  _RAND_135 = {1{`RANDOM}};
  way0Tag_6 = _RAND_135[20:0];
  _RAND_136 = {1{`RANDOM}};
  way0Tag_7 = _RAND_136[20:0];
  _RAND_137 = {1{`RANDOM}};
  way0Tag_8 = _RAND_137[20:0];
  _RAND_138 = {1{`RANDOM}};
  way0Tag_9 = _RAND_138[20:0];
  _RAND_139 = {1{`RANDOM}};
  way0Tag_10 = _RAND_139[20:0];
  _RAND_140 = {1{`RANDOM}};
  way0Tag_11 = _RAND_140[20:0];
  _RAND_141 = {1{`RANDOM}};
  way0Tag_12 = _RAND_141[20:0];
  _RAND_142 = {1{`RANDOM}};
  way0Tag_13 = _RAND_142[20:0];
  _RAND_143 = {1{`RANDOM}};
  way0Tag_14 = _RAND_143[20:0];
  _RAND_144 = {1{`RANDOM}};
  way0Tag_15 = _RAND_144[20:0];
  _RAND_145 = {1{`RANDOM}};
  way0Tag_16 = _RAND_145[20:0];
  _RAND_146 = {1{`RANDOM}};
  way0Tag_17 = _RAND_146[20:0];
  _RAND_147 = {1{`RANDOM}};
  way0Tag_18 = _RAND_147[20:0];
  _RAND_148 = {1{`RANDOM}};
  way0Tag_19 = _RAND_148[20:0];
  _RAND_149 = {1{`RANDOM}};
  way0Tag_20 = _RAND_149[20:0];
  _RAND_150 = {1{`RANDOM}};
  way0Tag_21 = _RAND_150[20:0];
  _RAND_151 = {1{`RANDOM}};
  way0Tag_22 = _RAND_151[20:0];
  _RAND_152 = {1{`RANDOM}};
  way0Tag_23 = _RAND_152[20:0];
  _RAND_153 = {1{`RANDOM}};
  way0Tag_24 = _RAND_153[20:0];
  _RAND_154 = {1{`RANDOM}};
  way0Tag_25 = _RAND_154[20:0];
  _RAND_155 = {1{`RANDOM}};
  way0Tag_26 = _RAND_155[20:0];
  _RAND_156 = {1{`RANDOM}};
  way0Tag_27 = _RAND_156[20:0];
  _RAND_157 = {1{`RANDOM}};
  way0Tag_28 = _RAND_157[20:0];
  _RAND_158 = {1{`RANDOM}};
  way0Tag_29 = _RAND_158[20:0];
  _RAND_159 = {1{`RANDOM}};
  way0Tag_30 = _RAND_159[20:0];
  _RAND_160 = {1{`RANDOM}};
  way0Tag_31 = _RAND_160[20:0];
  _RAND_161 = {1{`RANDOM}};
  way0Tag_32 = _RAND_161[20:0];
  _RAND_162 = {1{`RANDOM}};
  way0Tag_33 = _RAND_162[20:0];
  _RAND_163 = {1{`RANDOM}};
  way0Tag_34 = _RAND_163[20:0];
  _RAND_164 = {1{`RANDOM}};
  way0Tag_35 = _RAND_164[20:0];
  _RAND_165 = {1{`RANDOM}};
  way0Tag_36 = _RAND_165[20:0];
  _RAND_166 = {1{`RANDOM}};
  way0Tag_37 = _RAND_166[20:0];
  _RAND_167 = {1{`RANDOM}};
  way0Tag_38 = _RAND_167[20:0];
  _RAND_168 = {1{`RANDOM}};
  way0Tag_39 = _RAND_168[20:0];
  _RAND_169 = {1{`RANDOM}};
  way0Tag_40 = _RAND_169[20:0];
  _RAND_170 = {1{`RANDOM}};
  way0Tag_41 = _RAND_170[20:0];
  _RAND_171 = {1{`RANDOM}};
  way0Tag_42 = _RAND_171[20:0];
  _RAND_172 = {1{`RANDOM}};
  way0Tag_43 = _RAND_172[20:0];
  _RAND_173 = {1{`RANDOM}};
  way0Tag_44 = _RAND_173[20:0];
  _RAND_174 = {1{`RANDOM}};
  way0Tag_45 = _RAND_174[20:0];
  _RAND_175 = {1{`RANDOM}};
  way0Tag_46 = _RAND_175[20:0];
  _RAND_176 = {1{`RANDOM}};
  way0Tag_47 = _RAND_176[20:0];
  _RAND_177 = {1{`RANDOM}};
  way0Tag_48 = _RAND_177[20:0];
  _RAND_178 = {1{`RANDOM}};
  way0Tag_49 = _RAND_178[20:0];
  _RAND_179 = {1{`RANDOM}};
  way0Tag_50 = _RAND_179[20:0];
  _RAND_180 = {1{`RANDOM}};
  way0Tag_51 = _RAND_180[20:0];
  _RAND_181 = {1{`RANDOM}};
  way0Tag_52 = _RAND_181[20:0];
  _RAND_182 = {1{`RANDOM}};
  way0Tag_53 = _RAND_182[20:0];
  _RAND_183 = {1{`RANDOM}};
  way0Tag_54 = _RAND_183[20:0];
  _RAND_184 = {1{`RANDOM}};
  way0Tag_55 = _RAND_184[20:0];
  _RAND_185 = {1{`RANDOM}};
  way0Tag_56 = _RAND_185[20:0];
  _RAND_186 = {1{`RANDOM}};
  way0Tag_57 = _RAND_186[20:0];
  _RAND_187 = {1{`RANDOM}};
  way0Tag_58 = _RAND_187[20:0];
  _RAND_188 = {1{`RANDOM}};
  way0Tag_59 = _RAND_188[20:0];
  _RAND_189 = {1{`RANDOM}};
  way0Tag_60 = _RAND_189[20:0];
  _RAND_190 = {1{`RANDOM}};
  way0Tag_61 = _RAND_190[20:0];
  _RAND_191 = {1{`RANDOM}};
  way0Tag_62 = _RAND_191[20:0];
  _RAND_192 = {1{`RANDOM}};
  way0Tag_63 = _RAND_192[20:0];
  _RAND_193 = {1{`RANDOM}};
  way0Tag_64 = _RAND_193[20:0];
  _RAND_194 = {1{`RANDOM}};
  way0Tag_65 = _RAND_194[20:0];
  _RAND_195 = {1{`RANDOM}};
  way0Tag_66 = _RAND_195[20:0];
  _RAND_196 = {1{`RANDOM}};
  way0Tag_67 = _RAND_196[20:0];
  _RAND_197 = {1{`RANDOM}};
  way0Tag_68 = _RAND_197[20:0];
  _RAND_198 = {1{`RANDOM}};
  way0Tag_69 = _RAND_198[20:0];
  _RAND_199 = {1{`RANDOM}};
  way0Tag_70 = _RAND_199[20:0];
  _RAND_200 = {1{`RANDOM}};
  way0Tag_71 = _RAND_200[20:0];
  _RAND_201 = {1{`RANDOM}};
  way0Tag_72 = _RAND_201[20:0];
  _RAND_202 = {1{`RANDOM}};
  way0Tag_73 = _RAND_202[20:0];
  _RAND_203 = {1{`RANDOM}};
  way0Tag_74 = _RAND_203[20:0];
  _RAND_204 = {1{`RANDOM}};
  way0Tag_75 = _RAND_204[20:0];
  _RAND_205 = {1{`RANDOM}};
  way0Tag_76 = _RAND_205[20:0];
  _RAND_206 = {1{`RANDOM}};
  way0Tag_77 = _RAND_206[20:0];
  _RAND_207 = {1{`RANDOM}};
  way0Tag_78 = _RAND_207[20:0];
  _RAND_208 = {1{`RANDOM}};
  way0Tag_79 = _RAND_208[20:0];
  _RAND_209 = {1{`RANDOM}};
  way0Tag_80 = _RAND_209[20:0];
  _RAND_210 = {1{`RANDOM}};
  way0Tag_81 = _RAND_210[20:0];
  _RAND_211 = {1{`RANDOM}};
  way0Tag_82 = _RAND_211[20:0];
  _RAND_212 = {1{`RANDOM}};
  way0Tag_83 = _RAND_212[20:0];
  _RAND_213 = {1{`RANDOM}};
  way0Tag_84 = _RAND_213[20:0];
  _RAND_214 = {1{`RANDOM}};
  way0Tag_85 = _RAND_214[20:0];
  _RAND_215 = {1{`RANDOM}};
  way0Tag_86 = _RAND_215[20:0];
  _RAND_216 = {1{`RANDOM}};
  way0Tag_87 = _RAND_216[20:0];
  _RAND_217 = {1{`RANDOM}};
  way0Tag_88 = _RAND_217[20:0];
  _RAND_218 = {1{`RANDOM}};
  way0Tag_89 = _RAND_218[20:0];
  _RAND_219 = {1{`RANDOM}};
  way0Tag_90 = _RAND_219[20:0];
  _RAND_220 = {1{`RANDOM}};
  way0Tag_91 = _RAND_220[20:0];
  _RAND_221 = {1{`RANDOM}};
  way0Tag_92 = _RAND_221[20:0];
  _RAND_222 = {1{`RANDOM}};
  way0Tag_93 = _RAND_222[20:0];
  _RAND_223 = {1{`RANDOM}};
  way0Tag_94 = _RAND_223[20:0];
  _RAND_224 = {1{`RANDOM}};
  way0Tag_95 = _RAND_224[20:0];
  _RAND_225 = {1{`RANDOM}};
  way0Tag_96 = _RAND_225[20:0];
  _RAND_226 = {1{`RANDOM}};
  way0Tag_97 = _RAND_226[20:0];
  _RAND_227 = {1{`RANDOM}};
  way0Tag_98 = _RAND_227[20:0];
  _RAND_228 = {1{`RANDOM}};
  way0Tag_99 = _RAND_228[20:0];
  _RAND_229 = {1{`RANDOM}};
  way0Tag_100 = _RAND_229[20:0];
  _RAND_230 = {1{`RANDOM}};
  way0Tag_101 = _RAND_230[20:0];
  _RAND_231 = {1{`RANDOM}};
  way0Tag_102 = _RAND_231[20:0];
  _RAND_232 = {1{`RANDOM}};
  way0Tag_103 = _RAND_232[20:0];
  _RAND_233 = {1{`RANDOM}};
  way0Tag_104 = _RAND_233[20:0];
  _RAND_234 = {1{`RANDOM}};
  way0Tag_105 = _RAND_234[20:0];
  _RAND_235 = {1{`RANDOM}};
  way0Tag_106 = _RAND_235[20:0];
  _RAND_236 = {1{`RANDOM}};
  way0Tag_107 = _RAND_236[20:0];
  _RAND_237 = {1{`RANDOM}};
  way0Tag_108 = _RAND_237[20:0];
  _RAND_238 = {1{`RANDOM}};
  way0Tag_109 = _RAND_238[20:0];
  _RAND_239 = {1{`RANDOM}};
  way0Tag_110 = _RAND_239[20:0];
  _RAND_240 = {1{`RANDOM}};
  way0Tag_111 = _RAND_240[20:0];
  _RAND_241 = {1{`RANDOM}};
  way0Tag_112 = _RAND_241[20:0];
  _RAND_242 = {1{`RANDOM}};
  way0Tag_113 = _RAND_242[20:0];
  _RAND_243 = {1{`RANDOM}};
  way0Tag_114 = _RAND_243[20:0];
  _RAND_244 = {1{`RANDOM}};
  way0Tag_115 = _RAND_244[20:0];
  _RAND_245 = {1{`RANDOM}};
  way0Tag_116 = _RAND_245[20:0];
  _RAND_246 = {1{`RANDOM}};
  way0Tag_117 = _RAND_246[20:0];
  _RAND_247 = {1{`RANDOM}};
  way0Tag_118 = _RAND_247[20:0];
  _RAND_248 = {1{`RANDOM}};
  way0Tag_119 = _RAND_248[20:0];
  _RAND_249 = {1{`RANDOM}};
  way0Tag_120 = _RAND_249[20:0];
  _RAND_250 = {1{`RANDOM}};
  way0Tag_121 = _RAND_250[20:0];
  _RAND_251 = {1{`RANDOM}};
  way0Tag_122 = _RAND_251[20:0];
  _RAND_252 = {1{`RANDOM}};
  way0Tag_123 = _RAND_252[20:0];
  _RAND_253 = {1{`RANDOM}};
  way0Tag_124 = _RAND_253[20:0];
  _RAND_254 = {1{`RANDOM}};
  way0Tag_125 = _RAND_254[20:0];
  _RAND_255 = {1{`RANDOM}};
  way0Tag_126 = _RAND_255[20:0];
  _RAND_256 = {1{`RANDOM}};
  way0Tag_127 = _RAND_256[20:0];
  _RAND_257 = {1{`RANDOM}};
  way0Age_0 = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  way0Age_1 = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  way0Age_2 = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  way0Age_3 = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  way0Age_4 = _RAND_261[0:0];
  _RAND_262 = {1{`RANDOM}};
  way0Age_5 = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  way0Age_6 = _RAND_263[0:0];
  _RAND_264 = {1{`RANDOM}};
  way0Age_7 = _RAND_264[0:0];
  _RAND_265 = {1{`RANDOM}};
  way0Age_8 = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  way0Age_9 = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  way0Age_10 = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  way0Age_11 = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  way0Age_12 = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  way0Age_13 = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  way0Age_14 = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  way0Age_15 = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  way0Age_16 = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  way0Age_17 = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  way0Age_18 = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  way0Age_19 = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  way0Age_20 = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  way0Age_21 = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  way0Age_22 = _RAND_279[0:0];
  _RAND_280 = {1{`RANDOM}};
  way0Age_23 = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  way0Age_24 = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  way0Age_25 = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  way0Age_26 = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  way0Age_27 = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  way0Age_28 = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  way0Age_29 = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  way0Age_30 = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  way0Age_31 = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  way0Age_32 = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  way0Age_33 = _RAND_290[0:0];
  _RAND_291 = {1{`RANDOM}};
  way0Age_34 = _RAND_291[0:0];
  _RAND_292 = {1{`RANDOM}};
  way0Age_35 = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  way0Age_36 = _RAND_293[0:0];
  _RAND_294 = {1{`RANDOM}};
  way0Age_37 = _RAND_294[0:0];
  _RAND_295 = {1{`RANDOM}};
  way0Age_38 = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  way0Age_39 = _RAND_296[0:0];
  _RAND_297 = {1{`RANDOM}};
  way0Age_40 = _RAND_297[0:0];
  _RAND_298 = {1{`RANDOM}};
  way0Age_41 = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  way0Age_42 = _RAND_299[0:0];
  _RAND_300 = {1{`RANDOM}};
  way0Age_43 = _RAND_300[0:0];
  _RAND_301 = {1{`RANDOM}};
  way0Age_44 = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  way0Age_45 = _RAND_302[0:0];
  _RAND_303 = {1{`RANDOM}};
  way0Age_46 = _RAND_303[0:0];
  _RAND_304 = {1{`RANDOM}};
  way0Age_47 = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  way0Age_48 = _RAND_305[0:0];
  _RAND_306 = {1{`RANDOM}};
  way0Age_49 = _RAND_306[0:0];
  _RAND_307 = {1{`RANDOM}};
  way0Age_50 = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  way0Age_51 = _RAND_308[0:0];
  _RAND_309 = {1{`RANDOM}};
  way0Age_52 = _RAND_309[0:0];
  _RAND_310 = {1{`RANDOM}};
  way0Age_53 = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  way0Age_54 = _RAND_311[0:0];
  _RAND_312 = {1{`RANDOM}};
  way0Age_55 = _RAND_312[0:0];
  _RAND_313 = {1{`RANDOM}};
  way0Age_56 = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  way0Age_57 = _RAND_314[0:0];
  _RAND_315 = {1{`RANDOM}};
  way0Age_58 = _RAND_315[0:0];
  _RAND_316 = {1{`RANDOM}};
  way0Age_59 = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  way0Age_60 = _RAND_317[0:0];
  _RAND_318 = {1{`RANDOM}};
  way0Age_61 = _RAND_318[0:0];
  _RAND_319 = {1{`RANDOM}};
  way0Age_62 = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  way0Age_63 = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  way0Age_64 = _RAND_321[0:0];
  _RAND_322 = {1{`RANDOM}};
  way0Age_65 = _RAND_322[0:0];
  _RAND_323 = {1{`RANDOM}};
  way0Age_66 = _RAND_323[0:0];
  _RAND_324 = {1{`RANDOM}};
  way0Age_67 = _RAND_324[0:0];
  _RAND_325 = {1{`RANDOM}};
  way0Age_68 = _RAND_325[0:0];
  _RAND_326 = {1{`RANDOM}};
  way0Age_69 = _RAND_326[0:0];
  _RAND_327 = {1{`RANDOM}};
  way0Age_70 = _RAND_327[0:0];
  _RAND_328 = {1{`RANDOM}};
  way0Age_71 = _RAND_328[0:0];
  _RAND_329 = {1{`RANDOM}};
  way0Age_72 = _RAND_329[0:0];
  _RAND_330 = {1{`RANDOM}};
  way0Age_73 = _RAND_330[0:0];
  _RAND_331 = {1{`RANDOM}};
  way0Age_74 = _RAND_331[0:0];
  _RAND_332 = {1{`RANDOM}};
  way0Age_75 = _RAND_332[0:0];
  _RAND_333 = {1{`RANDOM}};
  way0Age_76 = _RAND_333[0:0];
  _RAND_334 = {1{`RANDOM}};
  way0Age_77 = _RAND_334[0:0];
  _RAND_335 = {1{`RANDOM}};
  way0Age_78 = _RAND_335[0:0];
  _RAND_336 = {1{`RANDOM}};
  way0Age_79 = _RAND_336[0:0];
  _RAND_337 = {1{`RANDOM}};
  way0Age_80 = _RAND_337[0:0];
  _RAND_338 = {1{`RANDOM}};
  way0Age_81 = _RAND_338[0:0];
  _RAND_339 = {1{`RANDOM}};
  way0Age_82 = _RAND_339[0:0];
  _RAND_340 = {1{`RANDOM}};
  way0Age_83 = _RAND_340[0:0];
  _RAND_341 = {1{`RANDOM}};
  way0Age_84 = _RAND_341[0:0];
  _RAND_342 = {1{`RANDOM}};
  way0Age_85 = _RAND_342[0:0];
  _RAND_343 = {1{`RANDOM}};
  way0Age_86 = _RAND_343[0:0];
  _RAND_344 = {1{`RANDOM}};
  way0Age_87 = _RAND_344[0:0];
  _RAND_345 = {1{`RANDOM}};
  way0Age_88 = _RAND_345[0:0];
  _RAND_346 = {1{`RANDOM}};
  way0Age_89 = _RAND_346[0:0];
  _RAND_347 = {1{`RANDOM}};
  way0Age_90 = _RAND_347[0:0];
  _RAND_348 = {1{`RANDOM}};
  way0Age_91 = _RAND_348[0:0];
  _RAND_349 = {1{`RANDOM}};
  way0Age_92 = _RAND_349[0:0];
  _RAND_350 = {1{`RANDOM}};
  way0Age_93 = _RAND_350[0:0];
  _RAND_351 = {1{`RANDOM}};
  way0Age_94 = _RAND_351[0:0];
  _RAND_352 = {1{`RANDOM}};
  way0Age_95 = _RAND_352[0:0];
  _RAND_353 = {1{`RANDOM}};
  way0Age_96 = _RAND_353[0:0];
  _RAND_354 = {1{`RANDOM}};
  way0Age_97 = _RAND_354[0:0];
  _RAND_355 = {1{`RANDOM}};
  way0Age_98 = _RAND_355[0:0];
  _RAND_356 = {1{`RANDOM}};
  way0Age_99 = _RAND_356[0:0];
  _RAND_357 = {1{`RANDOM}};
  way0Age_100 = _RAND_357[0:0];
  _RAND_358 = {1{`RANDOM}};
  way0Age_101 = _RAND_358[0:0];
  _RAND_359 = {1{`RANDOM}};
  way0Age_102 = _RAND_359[0:0];
  _RAND_360 = {1{`RANDOM}};
  way0Age_103 = _RAND_360[0:0];
  _RAND_361 = {1{`RANDOM}};
  way0Age_104 = _RAND_361[0:0];
  _RAND_362 = {1{`RANDOM}};
  way0Age_105 = _RAND_362[0:0];
  _RAND_363 = {1{`RANDOM}};
  way0Age_106 = _RAND_363[0:0];
  _RAND_364 = {1{`RANDOM}};
  way0Age_107 = _RAND_364[0:0];
  _RAND_365 = {1{`RANDOM}};
  way0Age_108 = _RAND_365[0:0];
  _RAND_366 = {1{`RANDOM}};
  way0Age_109 = _RAND_366[0:0];
  _RAND_367 = {1{`RANDOM}};
  way0Age_110 = _RAND_367[0:0];
  _RAND_368 = {1{`RANDOM}};
  way0Age_111 = _RAND_368[0:0];
  _RAND_369 = {1{`RANDOM}};
  way0Age_112 = _RAND_369[0:0];
  _RAND_370 = {1{`RANDOM}};
  way0Age_113 = _RAND_370[0:0];
  _RAND_371 = {1{`RANDOM}};
  way0Age_114 = _RAND_371[0:0];
  _RAND_372 = {1{`RANDOM}};
  way0Age_115 = _RAND_372[0:0];
  _RAND_373 = {1{`RANDOM}};
  way0Age_116 = _RAND_373[0:0];
  _RAND_374 = {1{`RANDOM}};
  way0Age_117 = _RAND_374[0:0];
  _RAND_375 = {1{`RANDOM}};
  way0Age_118 = _RAND_375[0:0];
  _RAND_376 = {1{`RANDOM}};
  way0Age_119 = _RAND_376[0:0];
  _RAND_377 = {1{`RANDOM}};
  way0Age_120 = _RAND_377[0:0];
  _RAND_378 = {1{`RANDOM}};
  way0Age_121 = _RAND_378[0:0];
  _RAND_379 = {1{`RANDOM}};
  way0Age_122 = _RAND_379[0:0];
  _RAND_380 = {1{`RANDOM}};
  way0Age_123 = _RAND_380[0:0];
  _RAND_381 = {1{`RANDOM}};
  way0Age_124 = _RAND_381[0:0];
  _RAND_382 = {1{`RANDOM}};
  way0Age_125 = _RAND_382[0:0];
  _RAND_383 = {1{`RANDOM}};
  way0Age_126 = _RAND_383[0:0];
  _RAND_384 = {1{`RANDOM}};
  way0Age_127 = _RAND_384[0:0];
  _RAND_385 = {1{`RANDOM}};
  way1V_0 = _RAND_385[0:0];
  _RAND_386 = {1{`RANDOM}};
  way1V_1 = _RAND_386[0:0];
  _RAND_387 = {1{`RANDOM}};
  way1V_2 = _RAND_387[0:0];
  _RAND_388 = {1{`RANDOM}};
  way1V_3 = _RAND_388[0:0];
  _RAND_389 = {1{`RANDOM}};
  way1V_4 = _RAND_389[0:0];
  _RAND_390 = {1{`RANDOM}};
  way1V_5 = _RAND_390[0:0];
  _RAND_391 = {1{`RANDOM}};
  way1V_6 = _RAND_391[0:0];
  _RAND_392 = {1{`RANDOM}};
  way1V_7 = _RAND_392[0:0];
  _RAND_393 = {1{`RANDOM}};
  way1V_8 = _RAND_393[0:0];
  _RAND_394 = {1{`RANDOM}};
  way1V_9 = _RAND_394[0:0];
  _RAND_395 = {1{`RANDOM}};
  way1V_10 = _RAND_395[0:0];
  _RAND_396 = {1{`RANDOM}};
  way1V_11 = _RAND_396[0:0];
  _RAND_397 = {1{`RANDOM}};
  way1V_12 = _RAND_397[0:0];
  _RAND_398 = {1{`RANDOM}};
  way1V_13 = _RAND_398[0:0];
  _RAND_399 = {1{`RANDOM}};
  way1V_14 = _RAND_399[0:0];
  _RAND_400 = {1{`RANDOM}};
  way1V_15 = _RAND_400[0:0];
  _RAND_401 = {1{`RANDOM}};
  way1V_16 = _RAND_401[0:0];
  _RAND_402 = {1{`RANDOM}};
  way1V_17 = _RAND_402[0:0];
  _RAND_403 = {1{`RANDOM}};
  way1V_18 = _RAND_403[0:0];
  _RAND_404 = {1{`RANDOM}};
  way1V_19 = _RAND_404[0:0];
  _RAND_405 = {1{`RANDOM}};
  way1V_20 = _RAND_405[0:0];
  _RAND_406 = {1{`RANDOM}};
  way1V_21 = _RAND_406[0:0];
  _RAND_407 = {1{`RANDOM}};
  way1V_22 = _RAND_407[0:0];
  _RAND_408 = {1{`RANDOM}};
  way1V_23 = _RAND_408[0:0];
  _RAND_409 = {1{`RANDOM}};
  way1V_24 = _RAND_409[0:0];
  _RAND_410 = {1{`RANDOM}};
  way1V_25 = _RAND_410[0:0];
  _RAND_411 = {1{`RANDOM}};
  way1V_26 = _RAND_411[0:0];
  _RAND_412 = {1{`RANDOM}};
  way1V_27 = _RAND_412[0:0];
  _RAND_413 = {1{`RANDOM}};
  way1V_28 = _RAND_413[0:0];
  _RAND_414 = {1{`RANDOM}};
  way1V_29 = _RAND_414[0:0];
  _RAND_415 = {1{`RANDOM}};
  way1V_30 = _RAND_415[0:0];
  _RAND_416 = {1{`RANDOM}};
  way1V_31 = _RAND_416[0:0];
  _RAND_417 = {1{`RANDOM}};
  way1V_32 = _RAND_417[0:0];
  _RAND_418 = {1{`RANDOM}};
  way1V_33 = _RAND_418[0:0];
  _RAND_419 = {1{`RANDOM}};
  way1V_34 = _RAND_419[0:0];
  _RAND_420 = {1{`RANDOM}};
  way1V_35 = _RAND_420[0:0];
  _RAND_421 = {1{`RANDOM}};
  way1V_36 = _RAND_421[0:0];
  _RAND_422 = {1{`RANDOM}};
  way1V_37 = _RAND_422[0:0];
  _RAND_423 = {1{`RANDOM}};
  way1V_38 = _RAND_423[0:0];
  _RAND_424 = {1{`RANDOM}};
  way1V_39 = _RAND_424[0:0];
  _RAND_425 = {1{`RANDOM}};
  way1V_40 = _RAND_425[0:0];
  _RAND_426 = {1{`RANDOM}};
  way1V_41 = _RAND_426[0:0];
  _RAND_427 = {1{`RANDOM}};
  way1V_42 = _RAND_427[0:0];
  _RAND_428 = {1{`RANDOM}};
  way1V_43 = _RAND_428[0:0];
  _RAND_429 = {1{`RANDOM}};
  way1V_44 = _RAND_429[0:0];
  _RAND_430 = {1{`RANDOM}};
  way1V_45 = _RAND_430[0:0];
  _RAND_431 = {1{`RANDOM}};
  way1V_46 = _RAND_431[0:0];
  _RAND_432 = {1{`RANDOM}};
  way1V_47 = _RAND_432[0:0];
  _RAND_433 = {1{`RANDOM}};
  way1V_48 = _RAND_433[0:0];
  _RAND_434 = {1{`RANDOM}};
  way1V_49 = _RAND_434[0:0];
  _RAND_435 = {1{`RANDOM}};
  way1V_50 = _RAND_435[0:0];
  _RAND_436 = {1{`RANDOM}};
  way1V_51 = _RAND_436[0:0];
  _RAND_437 = {1{`RANDOM}};
  way1V_52 = _RAND_437[0:0];
  _RAND_438 = {1{`RANDOM}};
  way1V_53 = _RAND_438[0:0];
  _RAND_439 = {1{`RANDOM}};
  way1V_54 = _RAND_439[0:0];
  _RAND_440 = {1{`RANDOM}};
  way1V_55 = _RAND_440[0:0];
  _RAND_441 = {1{`RANDOM}};
  way1V_56 = _RAND_441[0:0];
  _RAND_442 = {1{`RANDOM}};
  way1V_57 = _RAND_442[0:0];
  _RAND_443 = {1{`RANDOM}};
  way1V_58 = _RAND_443[0:0];
  _RAND_444 = {1{`RANDOM}};
  way1V_59 = _RAND_444[0:0];
  _RAND_445 = {1{`RANDOM}};
  way1V_60 = _RAND_445[0:0];
  _RAND_446 = {1{`RANDOM}};
  way1V_61 = _RAND_446[0:0];
  _RAND_447 = {1{`RANDOM}};
  way1V_62 = _RAND_447[0:0];
  _RAND_448 = {1{`RANDOM}};
  way1V_63 = _RAND_448[0:0];
  _RAND_449 = {1{`RANDOM}};
  way1V_64 = _RAND_449[0:0];
  _RAND_450 = {1{`RANDOM}};
  way1V_65 = _RAND_450[0:0];
  _RAND_451 = {1{`RANDOM}};
  way1V_66 = _RAND_451[0:0];
  _RAND_452 = {1{`RANDOM}};
  way1V_67 = _RAND_452[0:0];
  _RAND_453 = {1{`RANDOM}};
  way1V_68 = _RAND_453[0:0];
  _RAND_454 = {1{`RANDOM}};
  way1V_69 = _RAND_454[0:0];
  _RAND_455 = {1{`RANDOM}};
  way1V_70 = _RAND_455[0:0];
  _RAND_456 = {1{`RANDOM}};
  way1V_71 = _RAND_456[0:0];
  _RAND_457 = {1{`RANDOM}};
  way1V_72 = _RAND_457[0:0];
  _RAND_458 = {1{`RANDOM}};
  way1V_73 = _RAND_458[0:0];
  _RAND_459 = {1{`RANDOM}};
  way1V_74 = _RAND_459[0:0];
  _RAND_460 = {1{`RANDOM}};
  way1V_75 = _RAND_460[0:0];
  _RAND_461 = {1{`RANDOM}};
  way1V_76 = _RAND_461[0:0];
  _RAND_462 = {1{`RANDOM}};
  way1V_77 = _RAND_462[0:0];
  _RAND_463 = {1{`RANDOM}};
  way1V_78 = _RAND_463[0:0];
  _RAND_464 = {1{`RANDOM}};
  way1V_79 = _RAND_464[0:0];
  _RAND_465 = {1{`RANDOM}};
  way1V_80 = _RAND_465[0:0];
  _RAND_466 = {1{`RANDOM}};
  way1V_81 = _RAND_466[0:0];
  _RAND_467 = {1{`RANDOM}};
  way1V_82 = _RAND_467[0:0];
  _RAND_468 = {1{`RANDOM}};
  way1V_83 = _RAND_468[0:0];
  _RAND_469 = {1{`RANDOM}};
  way1V_84 = _RAND_469[0:0];
  _RAND_470 = {1{`RANDOM}};
  way1V_85 = _RAND_470[0:0];
  _RAND_471 = {1{`RANDOM}};
  way1V_86 = _RAND_471[0:0];
  _RAND_472 = {1{`RANDOM}};
  way1V_87 = _RAND_472[0:0];
  _RAND_473 = {1{`RANDOM}};
  way1V_88 = _RAND_473[0:0];
  _RAND_474 = {1{`RANDOM}};
  way1V_89 = _RAND_474[0:0];
  _RAND_475 = {1{`RANDOM}};
  way1V_90 = _RAND_475[0:0];
  _RAND_476 = {1{`RANDOM}};
  way1V_91 = _RAND_476[0:0];
  _RAND_477 = {1{`RANDOM}};
  way1V_92 = _RAND_477[0:0];
  _RAND_478 = {1{`RANDOM}};
  way1V_93 = _RAND_478[0:0];
  _RAND_479 = {1{`RANDOM}};
  way1V_94 = _RAND_479[0:0];
  _RAND_480 = {1{`RANDOM}};
  way1V_95 = _RAND_480[0:0];
  _RAND_481 = {1{`RANDOM}};
  way1V_96 = _RAND_481[0:0];
  _RAND_482 = {1{`RANDOM}};
  way1V_97 = _RAND_482[0:0];
  _RAND_483 = {1{`RANDOM}};
  way1V_98 = _RAND_483[0:0];
  _RAND_484 = {1{`RANDOM}};
  way1V_99 = _RAND_484[0:0];
  _RAND_485 = {1{`RANDOM}};
  way1V_100 = _RAND_485[0:0];
  _RAND_486 = {1{`RANDOM}};
  way1V_101 = _RAND_486[0:0];
  _RAND_487 = {1{`RANDOM}};
  way1V_102 = _RAND_487[0:0];
  _RAND_488 = {1{`RANDOM}};
  way1V_103 = _RAND_488[0:0];
  _RAND_489 = {1{`RANDOM}};
  way1V_104 = _RAND_489[0:0];
  _RAND_490 = {1{`RANDOM}};
  way1V_105 = _RAND_490[0:0];
  _RAND_491 = {1{`RANDOM}};
  way1V_106 = _RAND_491[0:0];
  _RAND_492 = {1{`RANDOM}};
  way1V_107 = _RAND_492[0:0];
  _RAND_493 = {1{`RANDOM}};
  way1V_108 = _RAND_493[0:0];
  _RAND_494 = {1{`RANDOM}};
  way1V_109 = _RAND_494[0:0];
  _RAND_495 = {1{`RANDOM}};
  way1V_110 = _RAND_495[0:0];
  _RAND_496 = {1{`RANDOM}};
  way1V_111 = _RAND_496[0:0];
  _RAND_497 = {1{`RANDOM}};
  way1V_112 = _RAND_497[0:0];
  _RAND_498 = {1{`RANDOM}};
  way1V_113 = _RAND_498[0:0];
  _RAND_499 = {1{`RANDOM}};
  way1V_114 = _RAND_499[0:0];
  _RAND_500 = {1{`RANDOM}};
  way1V_115 = _RAND_500[0:0];
  _RAND_501 = {1{`RANDOM}};
  way1V_116 = _RAND_501[0:0];
  _RAND_502 = {1{`RANDOM}};
  way1V_117 = _RAND_502[0:0];
  _RAND_503 = {1{`RANDOM}};
  way1V_118 = _RAND_503[0:0];
  _RAND_504 = {1{`RANDOM}};
  way1V_119 = _RAND_504[0:0];
  _RAND_505 = {1{`RANDOM}};
  way1V_120 = _RAND_505[0:0];
  _RAND_506 = {1{`RANDOM}};
  way1V_121 = _RAND_506[0:0];
  _RAND_507 = {1{`RANDOM}};
  way1V_122 = _RAND_507[0:0];
  _RAND_508 = {1{`RANDOM}};
  way1V_123 = _RAND_508[0:0];
  _RAND_509 = {1{`RANDOM}};
  way1V_124 = _RAND_509[0:0];
  _RAND_510 = {1{`RANDOM}};
  way1V_125 = _RAND_510[0:0];
  _RAND_511 = {1{`RANDOM}};
  way1V_126 = _RAND_511[0:0];
  _RAND_512 = {1{`RANDOM}};
  way1V_127 = _RAND_512[0:0];
  _RAND_513 = {1{`RANDOM}};
  way1Tag_0 = _RAND_513[20:0];
  _RAND_514 = {1{`RANDOM}};
  way1Tag_1 = _RAND_514[20:0];
  _RAND_515 = {1{`RANDOM}};
  way1Tag_2 = _RAND_515[20:0];
  _RAND_516 = {1{`RANDOM}};
  way1Tag_3 = _RAND_516[20:0];
  _RAND_517 = {1{`RANDOM}};
  way1Tag_4 = _RAND_517[20:0];
  _RAND_518 = {1{`RANDOM}};
  way1Tag_5 = _RAND_518[20:0];
  _RAND_519 = {1{`RANDOM}};
  way1Tag_6 = _RAND_519[20:0];
  _RAND_520 = {1{`RANDOM}};
  way1Tag_7 = _RAND_520[20:0];
  _RAND_521 = {1{`RANDOM}};
  way1Tag_8 = _RAND_521[20:0];
  _RAND_522 = {1{`RANDOM}};
  way1Tag_9 = _RAND_522[20:0];
  _RAND_523 = {1{`RANDOM}};
  way1Tag_10 = _RAND_523[20:0];
  _RAND_524 = {1{`RANDOM}};
  way1Tag_11 = _RAND_524[20:0];
  _RAND_525 = {1{`RANDOM}};
  way1Tag_12 = _RAND_525[20:0];
  _RAND_526 = {1{`RANDOM}};
  way1Tag_13 = _RAND_526[20:0];
  _RAND_527 = {1{`RANDOM}};
  way1Tag_14 = _RAND_527[20:0];
  _RAND_528 = {1{`RANDOM}};
  way1Tag_15 = _RAND_528[20:0];
  _RAND_529 = {1{`RANDOM}};
  way1Tag_16 = _RAND_529[20:0];
  _RAND_530 = {1{`RANDOM}};
  way1Tag_17 = _RAND_530[20:0];
  _RAND_531 = {1{`RANDOM}};
  way1Tag_18 = _RAND_531[20:0];
  _RAND_532 = {1{`RANDOM}};
  way1Tag_19 = _RAND_532[20:0];
  _RAND_533 = {1{`RANDOM}};
  way1Tag_20 = _RAND_533[20:0];
  _RAND_534 = {1{`RANDOM}};
  way1Tag_21 = _RAND_534[20:0];
  _RAND_535 = {1{`RANDOM}};
  way1Tag_22 = _RAND_535[20:0];
  _RAND_536 = {1{`RANDOM}};
  way1Tag_23 = _RAND_536[20:0];
  _RAND_537 = {1{`RANDOM}};
  way1Tag_24 = _RAND_537[20:0];
  _RAND_538 = {1{`RANDOM}};
  way1Tag_25 = _RAND_538[20:0];
  _RAND_539 = {1{`RANDOM}};
  way1Tag_26 = _RAND_539[20:0];
  _RAND_540 = {1{`RANDOM}};
  way1Tag_27 = _RAND_540[20:0];
  _RAND_541 = {1{`RANDOM}};
  way1Tag_28 = _RAND_541[20:0];
  _RAND_542 = {1{`RANDOM}};
  way1Tag_29 = _RAND_542[20:0];
  _RAND_543 = {1{`RANDOM}};
  way1Tag_30 = _RAND_543[20:0];
  _RAND_544 = {1{`RANDOM}};
  way1Tag_31 = _RAND_544[20:0];
  _RAND_545 = {1{`RANDOM}};
  way1Tag_32 = _RAND_545[20:0];
  _RAND_546 = {1{`RANDOM}};
  way1Tag_33 = _RAND_546[20:0];
  _RAND_547 = {1{`RANDOM}};
  way1Tag_34 = _RAND_547[20:0];
  _RAND_548 = {1{`RANDOM}};
  way1Tag_35 = _RAND_548[20:0];
  _RAND_549 = {1{`RANDOM}};
  way1Tag_36 = _RAND_549[20:0];
  _RAND_550 = {1{`RANDOM}};
  way1Tag_37 = _RAND_550[20:0];
  _RAND_551 = {1{`RANDOM}};
  way1Tag_38 = _RAND_551[20:0];
  _RAND_552 = {1{`RANDOM}};
  way1Tag_39 = _RAND_552[20:0];
  _RAND_553 = {1{`RANDOM}};
  way1Tag_40 = _RAND_553[20:0];
  _RAND_554 = {1{`RANDOM}};
  way1Tag_41 = _RAND_554[20:0];
  _RAND_555 = {1{`RANDOM}};
  way1Tag_42 = _RAND_555[20:0];
  _RAND_556 = {1{`RANDOM}};
  way1Tag_43 = _RAND_556[20:0];
  _RAND_557 = {1{`RANDOM}};
  way1Tag_44 = _RAND_557[20:0];
  _RAND_558 = {1{`RANDOM}};
  way1Tag_45 = _RAND_558[20:0];
  _RAND_559 = {1{`RANDOM}};
  way1Tag_46 = _RAND_559[20:0];
  _RAND_560 = {1{`RANDOM}};
  way1Tag_47 = _RAND_560[20:0];
  _RAND_561 = {1{`RANDOM}};
  way1Tag_48 = _RAND_561[20:0];
  _RAND_562 = {1{`RANDOM}};
  way1Tag_49 = _RAND_562[20:0];
  _RAND_563 = {1{`RANDOM}};
  way1Tag_50 = _RAND_563[20:0];
  _RAND_564 = {1{`RANDOM}};
  way1Tag_51 = _RAND_564[20:0];
  _RAND_565 = {1{`RANDOM}};
  way1Tag_52 = _RAND_565[20:0];
  _RAND_566 = {1{`RANDOM}};
  way1Tag_53 = _RAND_566[20:0];
  _RAND_567 = {1{`RANDOM}};
  way1Tag_54 = _RAND_567[20:0];
  _RAND_568 = {1{`RANDOM}};
  way1Tag_55 = _RAND_568[20:0];
  _RAND_569 = {1{`RANDOM}};
  way1Tag_56 = _RAND_569[20:0];
  _RAND_570 = {1{`RANDOM}};
  way1Tag_57 = _RAND_570[20:0];
  _RAND_571 = {1{`RANDOM}};
  way1Tag_58 = _RAND_571[20:0];
  _RAND_572 = {1{`RANDOM}};
  way1Tag_59 = _RAND_572[20:0];
  _RAND_573 = {1{`RANDOM}};
  way1Tag_60 = _RAND_573[20:0];
  _RAND_574 = {1{`RANDOM}};
  way1Tag_61 = _RAND_574[20:0];
  _RAND_575 = {1{`RANDOM}};
  way1Tag_62 = _RAND_575[20:0];
  _RAND_576 = {1{`RANDOM}};
  way1Tag_63 = _RAND_576[20:0];
  _RAND_577 = {1{`RANDOM}};
  way1Tag_64 = _RAND_577[20:0];
  _RAND_578 = {1{`RANDOM}};
  way1Tag_65 = _RAND_578[20:0];
  _RAND_579 = {1{`RANDOM}};
  way1Tag_66 = _RAND_579[20:0];
  _RAND_580 = {1{`RANDOM}};
  way1Tag_67 = _RAND_580[20:0];
  _RAND_581 = {1{`RANDOM}};
  way1Tag_68 = _RAND_581[20:0];
  _RAND_582 = {1{`RANDOM}};
  way1Tag_69 = _RAND_582[20:0];
  _RAND_583 = {1{`RANDOM}};
  way1Tag_70 = _RAND_583[20:0];
  _RAND_584 = {1{`RANDOM}};
  way1Tag_71 = _RAND_584[20:0];
  _RAND_585 = {1{`RANDOM}};
  way1Tag_72 = _RAND_585[20:0];
  _RAND_586 = {1{`RANDOM}};
  way1Tag_73 = _RAND_586[20:0];
  _RAND_587 = {1{`RANDOM}};
  way1Tag_74 = _RAND_587[20:0];
  _RAND_588 = {1{`RANDOM}};
  way1Tag_75 = _RAND_588[20:0];
  _RAND_589 = {1{`RANDOM}};
  way1Tag_76 = _RAND_589[20:0];
  _RAND_590 = {1{`RANDOM}};
  way1Tag_77 = _RAND_590[20:0];
  _RAND_591 = {1{`RANDOM}};
  way1Tag_78 = _RAND_591[20:0];
  _RAND_592 = {1{`RANDOM}};
  way1Tag_79 = _RAND_592[20:0];
  _RAND_593 = {1{`RANDOM}};
  way1Tag_80 = _RAND_593[20:0];
  _RAND_594 = {1{`RANDOM}};
  way1Tag_81 = _RAND_594[20:0];
  _RAND_595 = {1{`RANDOM}};
  way1Tag_82 = _RAND_595[20:0];
  _RAND_596 = {1{`RANDOM}};
  way1Tag_83 = _RAND_596[20:0];
  _RAND_597 = {1{`RANDOM}};
  way1Tag_84 = _RAND_597[20:0];
  _RAND_598 = {1{`RANDOM}};
  way1Tag_85 = _RAND_598[20:0];
  _RAND_599 = {1{`RANDOM}};
  way1Tag_86 = _RAND_599[20:0];
  _RAND_600 = {1{`RANDOM}};
  way1Tag_87 = _RAND_600[20:0];
  _RAND_601 = {1{`RANDOM}};
  way1Tag_88 = _RAND_601[20:0];
  _RAND_602 = {1{`RANDOM}};
  way1Tag_89 = _RAND_602[20:0];
  _RAND_603 = {1{`RANDOM}};
  way1Tag_90 = _RAND_603[20:0];
  _RAND_604 = {1{`RANDOM}};
  way1Tag_91 = _RAND_604[20:0];
  _RAND_605 = {1{`RANDOM}};
  way1Tag_92 = _RAND_605[20:0];
  _RAND_606 = {1{`RANDOM}};
  way1Tag_93 = _RAND_606[20:0];
  _RAND_607 = {1{`RANDOM}};
  way1Tag_94 = _RAND_607[20:0];
  _RAND_608 = {1{`RANDOM}};
  way1Tag_95 = _RAND_608[20:0];
  _RAND_609 = {1{`RANDOM}};
  way1Tag_96 = _RAND_609[20:0];
  _RAND_610 = {1{`RANDOM}};
  way1Tag_97 = _RAND_610[20:0];
  _RAND_611 = {1{`RANDOM}};
  way1Tag_98 = _RAND_611[20:0];
  _RAND_612 = {1{`RANDOM}};
  way1Tag_99 = _RAND_612[20:0];
  _RAND_613 = {1{`RANDOM}};
  way1Tag_100 = _RAND_613[20:0];
  _RAND_614 = {1{`RANDOM}};
  way1Tag_101 = _RAND_614[20:0];
  _RAND_615 = {1{`RANDOM}};
  way1Tag_102 = _RAND_615[20:0];
  _RAND_616 = {1{`RANDOM}};
  way1Tag_103 = _RAND_616[20:0];
  _RAND_617 = {1{`RANDOM}};
  way1Tag_104 = _RAND_617[20:0];
  _RAND_618 = {1{`RANDOM}};
  way1Tag_105 = _RAND_618[20:0];
  _RAND_619 = {1{`RANDOM}};
  way1Tag_106 = _RAND_619[20:0];
  _RAND_620 = {1{`RANDOM}};
  way1Tag_107 = _RAND_620[20:0];
  _RAND_621 = {1{`RANDOM}};
  way1Tag_108 = _RAND_621[20:0];
  _RAND_622 = {1{`RANDOM}};
  way1Tag_109 = _RAND_622[20:0];
  _RAND_623 = {1{`RANDOM}};
  way1Tag_110 = _RAND_623[20:0];
  _RAND_624 = {1{`RANDOM}};
  way1Tag_111 = _RAND_624[20:0];
  _RAND_625 = {1{`RANDOM}};
  way1Tag_112 = _RAND_625[20:0];
  _RAND_626 = {1{`RANDOM}};
  way1Tag_113 = _RAND_626[20:0];
  _RAND_627 = {1{`RANDOM}};
  way1Tag_114 = _RAND_627[20:0];
  _RAND_628 = {1{`RANDOM}};
  way1Tag_115 = _RAND_628[20:0];
  _RAND_629 = {1{`RANDOM}};
  way1Tag_116 = _RAND_629[20:0];
  _RAND_630 = {1{`RANDOM}};
  way1Tag_117 = _RAND_630[20:0];
  _RAND_631 = {1{`RANDOM}};
  way1Tag_118 = _RAND_631[20:0];
  _RAND_632 = {1{`RANDOM}};
  way1Tag_119 = _RAND_632[20:0];
  _RAND_633 = {1{`RANDOM}};
  way1Tag_120 = _RAND_633[20:0];
  _RAND_634 = {1{`RANDOM}};
  way1Tag_121 = _RAND_634[20:0];
  _RAND_635 = {1{`RANDOM}};
  way1Tag_122 = _RAND_635[20:0];
  _RAND_636 = {1{`RANDOM}};
  way1Tag_123 = _RAND_636[20:0];
  _RAND_637 = {1{`RANDOM}};
  way1Tag_124 = _RAND_637[20:0];
  _RAND_638 = {1{`RANDOM}};
  way1Tag_125 = _RAND_638[20:0];
  _RAND_639 = {1{`RANDOM}};
  way1Tag_126 = _RAND_639[20:0];
  _RAND_640 = {1{`RANDOM}};
  way1Tag_127 = _RAND_640[20:0];
  _RAND_641 = {1{`RANDOM}};
  way1Age_0 = _RAND_641[0:0];
  _RAND_642 = {1{`RANDOM}};
  way1Age_1 = _RAND_642[0:0];
  _RAND_643 = {1{`RANDOM}};
  way1Age_2 = _RAND_643[0:0];
  _RAND_644 = {1{`RANDOM}};
  way1Age_3 = _RAND_644[0:0];
  _RAND_645 = {1{`RANDOM}};
  way1Age_4 = _RAND_645[0:0];
  _RAND_646 = {1{`RANDOM}};
  way1Age_5 = _RAND_646[0:0];
  _RAND_647 = {1{`RANDOM}};
  way1Age_6 = _RAND_647[0:0];
  _RAND_648 = {1{`RANDOM}};
  way1Age_7 = _RAND_648[0:0];
  _RAND_649 = {1{`RANDOM}};
  way1Age_8 = _RAND_649[0:0];
  _RAND_650 = {1{`RANDOM}};
  way1Age_9 = _RAND_650[0:0];
  _RAND_651 = {1{`RANDOM}};
  way1Age_10 = _RAND_651[0:0];
  _RAND_652 = {1{`RANDOM}};
  way1Age_11 = _RAND_652[0:0];
  _RAND_653 = {1{`RANDOM}};
  way1Age_12 = _RAND_653[0:0];
  _RAND_654 = {1{`RANDOM}};
  way1Age_13 = _RAND_654[0:0];
  _RAND_655 = {1{`RANDOM}};
  way1Age_14 = _RAND_655[0:0];
  _RAND_656 = {1{`RANDOM}};
  way1Age_15 = _RAND_656[0:0];
  _RAND_657 = {1{`RANDOM}};
  way1Age_16 = _RAND_657[0:0];
  _RAND_658 = {1{`RANDOM}};
  way1Age_17 = _RAND_658[0:0];
  _RAND_659 = {1{`RANDOM}};
  way1Age_18 = _RAND_659[0:0];
  _RAND_660 = {1{`RANDOM}};
  way1Age_19 = _RAND_660[0:0];
  _RAND_661 = {1{`RANDOM}};
  way1Age_20 = _RAND_661[0:0];
  _RAND_662 = {1{`RANDOM}};
  way1Age_21 = _RAND_662[0:0];
  _RAND_663 = {1{`RANDOM}};
  way1Age_22 = _RAND_663[0:0];
  _RAND_664 = {1{`RANDOM}};
  way1Age_23 = _RAND_664[0:0];
  _RAND_665 = {1{`RANDOM}};
  way1Age_24 = _RAND_665[0:0];
  _RAND_666 = {1{`RANDOM}};
  way1Age_25 = _RAND_666[0:0];
  _RAND_667 = {1{`RANDOM}};
  way1Age_26 = _RAND_667[0:0];
  _RAND_668 = {1{`RANDOM}};
  way1Age_27 = _RAND_668[0:0];
  _RAND_669 = {1{`RANDOM}};
  way1Age_28 = _RAND_669[0:0];
  _RAND_670 = {1{`RANDOM}};
  way1Age_29 = _RAND_670[0:0];
  _RAND_671 = {1{`RANDOM}};
  way1Age_30 = _RAND_671[0:0];
  _RAND_672 = {1{`RANDOM}};
  way1Age_31 = _RAND_672[0:0];
  _RAND_673 = {1{`RANDOM}};
  way1Age_32 = _RAND_673[0:0];
  _RAND_674 = {1{`RANDOM}};
  way1Age_33 = _RAND_674[0:0];
  _RAND_675 = {1{`RANDOM}};
  way1Age_34 = _RAND_675[0:0];
  _RAND_676 = {1{`RANDOM}};
  way1Age_35 = _RAND_676[0:0];
  _RAND_677 = {1{`RANDOM}};
  way1Age_36 = _RAND_677[0:0];
  _RAND_678 = {1{`RANDOM}};
  way1Age_37 = _RAND_678[0:0];
  _RAND_679 = {1{`RANDOM}};
  way1Age_38 = _RAND_679[0:0];
  _RAND_680 = {1{`RANDOM}};
  way1Age_39 = _RAND_680[0:0];
  _RAND_681 = {1{`RANDOM}};
  way1Age_40 = _RAND_681[0:0];
  _RAND_682 = {1{`RANDOM}};
  way1Age_41 = _RAND_682[0:0];
  _RAND_683 = {1{`RANDOM}};
  way1Age_42 = _RAND_683[0:0];
  _RAND_684 = {1{`RANDOM}};
  way1Age_43 = _RAND_684[0:0];
  _RAND_685 = {1{`RANDOM}};
  way1Age_44 = _RAND_685[0:0];
  _RAND_686 = {1{`RANDOM}};
  way1Age_45 = _RAND_686[0:0];
  _RAND_687 = {1{`RANDOM}};
  way1Age_46 = _RAND_687[0:0];
  _RAND_688 = {1{`RANDOM}};
  way1Age_47 = _RAND_688[0:0];
  _RAND_689 = {1{`RANDOM}};
  way1Age_48 = _RAND_689[0:0];
  _RAND_690 = {1{`RANDOM}};
  way1Age_49 = _RAND_690[0:0];
  _RAND_691 = {1{`RANDOM}};
  way1Age_50 = _RAND_691[0:0];
  _RAND_692 = {1{`RANDOM}};
  way1Age_51 = _RAND_692[0:0];
  _RAND_693 = {1{`RANDOM}};
  way1Age_52 = _RAND_693[0:0];
  _RAND_694 = {1{`RANDOM}};
  way1Age_53 = _RAND_694[0:0];
  _RAND_695 = {1{`RANDOM}};
  way1Age_54 = _RAND_695[0:0];
  _RAND_696 = {1{`RANDOM}};
  way1Age_55 = _RAND_696[0:0];
  _RAND_697 = {1{`RANDOM}};
  way1Age_56 = _RAND_697[0:0];
  _RAND_698 = {1{`RANDOM}};
  way1Age_57 = _RAND_698[0:0];
  _RAND_699 = {1{`RANDOM}};
  way1Age_58 = _RAND_699[0:0];
  _RAND_700 = {1{`RANDOM}};
  way1Age_59 = _RAND_700[0:0];
  _RAND_701 = {1{`RANDOM}};
  way1Age_60 = _RAND_701[0:0];
  _RAND_702 = {1{`RANDOM}};
  way1Age_61 = _RAND_702[0:0];
  _RAND_703 = {1{`RANDOM}};
  way1Age_62 = _RAND_703[0:0];
  _RAND_704 = {1{`RANDOM}};
  way1Age_63 = _RAND_704[0:0];
  _RAND_705 = {1{`RANDOM}};
  way1Age_64 = _RAND_705[0:0];
  _RAND_706 = {1{`RANDOM}};
  way1Age_65 = _RAND_706[0:0];
  _RAND_707 = {1{`RANDOM}};
  way1Age_66 = _RAND_707[0:0];
  _RAND_708 = {1{`RANDOM}};
  way1Age_67 = _RAND_708[0:0];
  _RAND_709 = {1{`RANDOM}};
  way1Age_68 = _RAND_709[0:0];
  _RAND_710 = {1{`RANDOM}};
  way1Age_69 = _RAND_710[0:0];
  _RAND_711 = {1{`RANDOM}};
  way1Age_70 = _RAND_711[0:0];
  _RAND_712 = {1{`RANDOM}};
  way1Age_71 = _RAND_712[0:0];
  _RAND_713 = {1{`RANDOM}};
  way1Age_72 = _RAND_713[0:0];
  _RAND_714 = {1{`RANDOM}};
  way1Age_73 = _RAND_714[0:0];
  _RAND_715 = {1{`RANDOM}};
  way1Age_74 = _RAND_715[0:0];
  _RAND_716 = {1{`RANDOM}};
  way1Age_75 = _RAND_716[0:0];
  _RAND_717 = {1{`RANDOM}};
  way1Age_76 = _RAND_717[0:0];
  _RAND_718 = {1{`RANDOM}};
  way1Age_77 = _RAND_718[0:0];
  _RAND_719 = {1{`RANDOM}};
  way1Age_78 = _RAND_719[0:0];
  _RAND_720 = {1{`RANDOM}};
  way1Age_79 = _RAND_720[0:0];
  _RAND_721 = {1{`RANDOM}};
  way1Age_80 = _RAND_721[0:0];
  _RAND_722 = {1{`RANDOM}};
  way1Age_81 = _RAND_722[0:0];
  _RAND_723 = {1{`RANDOM}};
  way1Age_82 = _RAND_723[0:0];
  _RAND_724 = {1{`RANDOM}};
  way1Age_83 = _RAND_724[0:0];
  _RAND_725 = {1{`RANDOM}};
  way1Age_84 = _RAND_725[0:0];
  _RAND_726 = {1{`RANDOM}};
  way1Age_85 = _RAND_726[0:0];
  _RAND_727 = {1{`RANDOM}};
  way1Age_86 = _RAND_727[0:0];
  _RAND_728 = {1{`RANDOM}};
  way1Age_87 = _RAND_728[0:0];
  _RAND_729 = {1{`RANDOM}};
  way1Age_88 = _RAND_729[0:0];
  _RAND_730 = {1{`RANDOM}};
  way1Age_89 = _RAND_730[0:0];
  _RAND_731 = {1{`RANDOM}};
  way1Age_90 = _RAND_731[0:0];
  _RAND_732 = {1{`RANDOM}};
  way1Age_91 = _RAND_732[0:0];
  _RAND_733 = {1{`RANDOM}};
  way1Age_92 = _RAND_733[0:0];
  _RAND_734 = {1{`RANDOM}};
  way1Age_93 = _RAND_734[0:0];
  _RAND_735 = {1{`RANDOM}};
  way1Age_94 = _RAND_735[0:0];
  _RAND_736 = {1{`RANDOM}};
  way1Age_95 = _RAND_736[0:0];
  _RAND_737 = {1{`RANDOM}};
  way1Age_96 = _RAND_737[0:0];
  _RAND_738 = {1{`RANDOM}};
  way1Age_97 = _RAND_738[0:0];
  _RAND_739 = {1{`RANDOM}};
  way1Age_98 = _RAND_739[0:0];
  _RAND_740 = {1{`RANDOM}};
  way1Age_99 = _RAND_740[0:0];
  _RAND_741 = {1{`RANDOM}};
  way1Age_100 = _RAND_741[0:0];
  _RAND_742 = {1{`RANDOM}};
  way1Age_101 = _RAND_742[0:0];
  _RAND_743 = {1{`RANDOM}};
  way1Age_102 = _RAND_743[0:0];
  _RAND_744 = {1{`RANDOM}};
  way1Age_103 = _RAND_744[0:0];
  _RAND_745 = {1{`RANDOM}};
  way1Age_104 = _RAND_745[0:0];
  _RAND_746 = {1{`RANDOM}};
  way1Age_105 = _RAND_746[0:0];
  _RAND_747 = {1{`RANDOM}};
  way1Age_106 = _RAND_747[0:0];
  _RAND_748 = {1{`RANDOM}};
  way1Age_107 = _RAND_748[0:0];
  _RAND_749 = {1{`RANDOM}};
  way1Age_108 = _RAND_749[0:0];
  _RAND_750 = {1{`RANDOM}};
  way1Age_109 = _RAND_750[0:0];
  _RAND_751 = {1{`RANDOM}};
  way1Age_110 = _RAND_751[0:0];
  _RAND_752 = {1{`RANDOM}};
  way1Age_111 = _RAND_752[0:0];
  _RAND_753 = {1{`RANDOM}};
  way1Age_112 = _RAND_753[0:0];
  _RAND_754 = {1{`RANDOM}};
  way1Age_113 = _RAND_754[0:0];
  _RAND_755 = {1{`RANDOM}};
  way1Age_114 = _RAND_755[0:0];
  _RAND_756 = {1{`RANDOM}};
  way1Age_115 = _RAND_756[0:0];
  _RAND_757 = {1{`RANDOM}};
  way1Age_116 = _RAND_757[0:0];
  _RAND_758 = {1{`RANDOM}};
  way1Age_117 = _RAND_758[0:0];
  _RAND_759 = {1{`RANDOM}};
  way1Age_118 = _RAND_759[0:0];
  _RAND_760 = {1{`RANDOM}};
  way1Age_119 = _RAND_760[0:0];
  _RAND_761 = {1{`RANDOM}};
  way1Age_120 = _RAND_761[0:0];
  _RAND_762 = {1{`RANDOM}};
  way1Age_121 = _RAND_762[0:0];
  _RAND_763 = {1{`RANDOM}};
  way1Age_122 = _RAND_763[0:0];
  _RAND_764 = {1{`RANDOM}};
  way1Age_123 = _RAND_764[0:0];
  _RAND_765 = {1{`RANDOM}};
  way1Age_124 = _RAND_765[0:0];
  _RAND_766 = {1{`RANDOM}};
  way1Age_125 = _RAND_766[0:0];
  _RAND_767 = {1{`RANDOM}};
  way1Age_126 = _RAND_767[0:0];
  _RAND_768 = {1{`RANDOM}};
  way1Age_127 = _RAND_768[0:0];
  _RAND_769 = {1{`RANDOM}};
  state = _RAND_769[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module DCache(
  input          clock,
  input          reset,
  input          io_dmem_data_valid,
  output         io_dmem_data_ready,
  input          io_dmem_data_req,
  input  [31:0]  io_dmem_data_addr,
  input  [1:0]   io_dmem_data_size,
  input  [7:0]   io_dmem_data_strb,
  output [63:0]  io_dmem_data_read,
  input  [127:0] io_dmem_data_write,
  output         io_out_data_valid,
  input          io_out_data_ready,
  output         io_out_data_req,
  output [31:0]  io_out_data_addr,
  output [7:0]   io_out_data_strb,
  input  [127:0] io_out_data_read,
  output [127:0] io_out_data_write
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_645;
  reg [31:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_649;
  reg [31:0] _RAND_650;
  reg [31:0] _RAND_651;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
  reg [31:0] _RAND_654;
  reg [31:0] _RAND_655;
  reg [31:0] _RAND_656;
  reg [31:0] _RAND_657;
  reg [31:0] _RAND_658;
  reg [31:0] _RAND_659;
  reg [31:0] _RAND_660;
  reg [31:0] _RAND_661;
  reg [31:0] _RAND_662;
  reg [31:0] _RAND_663;
  reg [31:0] _RAND_664;
  reg [31:0] _RAND_665;
  reg [31:0] _RAND_666;
  reg [31:0] _RAND_667;
  reg [31:0] _RAND_668;
  reg [31:0] _RAND_669;
  reg [31:0] _RAND_670;
  reg [31:0] _RAND_671;
  reg [31:0] _RAND_672;
  reg [31:0] _RAND_673;
  reg [31:0] _RAND_674;
  reg [31:0] _RAND_675;
  reg [31:0] _RAND_676;
  reg [31:0] _RAND_677;
  reg [31:0] _RAND_678;
  reg [31:0] _RAND_679;
  reg [31:0] _RAND_680;
  reg [31:0] _RAND_681;
  reg [31:0] _RAND_682;
  reg [31:0] _RAND_683;
  reg [31:0] _RAND_684;
  reg [31:0] _RAND_685;
  reg [31:0] _RAND_686;
  reg [31:0] _RAND_687;
  reg [31:0] _RAND_688;
  reg [31:0] _RAND_689;
  reg [31:0] _RAND_690;
  reg [31:0] _RAND_691;
  reg [31:0] _RAND_692;
  reg [31:0] _RAND_693;
  reg [31:0] _RAND_694;
  reg [31:0] _RAND_695;
  reg [31:0] _RAND_696;
  reg [31:0] _RAND_697;
  reg [31:0] _RAND_698;
  reg [31:0] _RAND_699;
  reg [31:0] _RAND_700;
  reg [31:0] _RAND_701;
  reg [31:0] _RAND_702;
  reg [31:0] _RAND_703;
  reg [31:0] _RAND_704;
  reg [31:0] _RAND_705;
  reg [31:0] _RAND_706;
  reg [31:0] _RAND_707;
  reg [31:0] _RAND_708;
  reg [31:0] _RAND_709;
  reg [31:0] _RAND_710;
  reg [31:0] _RAND_711;
  reg [31:0] _RAND_712;
  reg [31:0] _RAND_713;
  reg [31:0] _RAND_714;
  reg [31:0] _RAND_715;
  reg [31:0] _RAND_716;
  reg [31:0] _RAND_717;
  reg [31:0] _RAND_718;
  reg [31:0] _RAND_719;
  reg [31:0] _RAND_720;
  reg [31:0] _RAND_721;
  reg [31:0] _RAND_722;
  reg [31:0] _RAND_723;
  reg [31:0] _RAND_724;
  reg [31:0] _RAND_725;
  reg [31:0] _RAND_726;
  reg [31:0] _RAND_727;
  reg [31:0] _RAND_728;
  reg [31:0] _RAND_729;
  reg [31:0] _RAND_730;
  reg [31:0] _RAND_731;
  reg [31:0] _RAND_732;
  reg [31:0] _RAND_733;
  reg [31:0] _RAND_734;
  reg [31:0] _RAND_735;
  reg [31:0] _RAND_736;
  reg [31:0] _RAND_737;
  reg [31:0] _RAND_738;
  reg [31:0] _RAND_739;
  reg [31:0] _RAND_740;
  reg [31:0] _RAND_741;
  reg [31:0] _RAND_742;
  reg [31:0] _RAND_743;
  reg [31:0] _RAND_744;
  reg [31:0] _RAND_745;
  reg [31:0] _RAND_746;
  reg [31:0] _RAND_747;
  reg [31:0] _RAND_748;
  reg [31:0] _RAND_749;
  reg [31:0] _RAND_750;
  reg [31:0] _RAND_751;
  reg [31:0] _RAND_752;
  reg [31:0] _RAND_753;
  reg [31:0] _RAND_754;
  reg [31:0] _RAND_755;
  reg [31:0] _RAND_756;
  reg [31:0] _RAND_757;
  reg [31:0] _RAND_758;
  reg [31:0] _RAND_759;
  reg [31:0] _RAND_760;
  reg [31:0] _RAND_761;
  reg [31:0] _RAND_762;
  reg [31:0] _RAND_763;
  reg [31:0] _RAND_764;
  reg [31:0] _RAND_765;
  reg [31:0] _RAND_766;
  reg [31:0] _RAND_767;
  reg [31:0] _RAND_768;
  reg [31:0] _RAND_769;
  reg [31:0] _RAND_770;
  reg [31:0] _RAND_771;
  reg [31:0] _RAND_772;
  reg [31:0] _RAND_773;
  reg [31:0] _RAND_774;
  reg [31:0] _RAND_775;
  reg [31:0] _RAND_776;
  reg [31:0] _RAND_777;
  reg [31:0] _RAND_778;
  reg [31:0] _RAND_779;
  reg [31:0] _RAND_780;
  reg [31:0] _RAND_781;
  reg [31:0] _RAND_782;
  reg [31:0] _RAND_783;
  reg [31:0] _RAND_784;
  reg [31:0] _RAND_785;
  reg [31:0] _RAND_786;
  reg [31:0] _RAND_787;
  reg [31:0] _RAND_788;
  reg [31:0] _RAND_789;
  reg [31:0] _RAND_790;
  reg [31:0] _RAND_791;
  reg [31:0] _RAND_792;
  reg [31:0] _RAND_793;
  reg [31:0] _RAND_794;
  reg [31:0] _RAND_795;
  reg [31:0] _RAND_796;
  reg [31:0] _RAND_797;
  reg [31:0] _RAND_798;
  reg [31:0] _RAND_799;
  reg [31:0] _RAND_800;
  reg [31:0] _RAND_801;
  reg [31:0] _RAND_802;
  reg [31:0] _RAND_803;
  reg [31:0] _RAND_804;
  reg [31:0] _RAND_805;
  reg [31:0] _RAND_806;
  reg [31:0] _RAND_807;
  reg [31:0] _RAND_808;
  reg [31:0] _RAND_809;
  reg [31:0] _RAND_810;
  reg [31:0] _RAND_811;
  reg [31:0] _RAND_812;
  reg [31:0] _RAND_813;
  reg [31:0] _RAND_814;
  reg [31:0] _RAND_815;
  reg [31:0] _RAND_816;
  reg [31:0] _RAND_817;
  reg [31:0] _RAND_818;
  reg [31:0] _RAND_819;
  reg [31:0] _RAND_820;
  reg [31:0] _RAND_821;
  reg [31:0] _RAND_822;
  reg [31:0] _RAND_823;
  reg [31:0] _RAND_824;
  reg [31:0] _RAND_825;
  reg [31:0] _RAND_826;
  reg [31:0] _RAND_827;
  reg [31:0] _RAND_828;
  reg [31:0] _RAND_829;
  reg [31:0] _RAND_830;
  reg [31:0] _RAND_831;
  reg [31:0] _RAND_832;
  reg [31:0] _RAND_833;
  reg [31:0] _RAND_834;
  reg [31:0] _RAND_835;
  reg [31:0] _RAND_836;
  reg [31:0] _RAND_837;
  reg [31:0] _RAND_838;
  reg [31:0] _RAND_839;
  reg [31:0] _RAND_840;
  reg [31:0] _RAND_841;
  reg [31:0] _RAND_842;
  reg [31:0] _RAND_843;
  reg [31:0] _RAND_844;
  reg [31:0] _RAND_845;
  reg [31:0] _RAND_846;
  reg [31:0] _RAND_847;
  reg [31:0] _RAND_848;
  reg [31:0] _RAND_849;
  reg [31:0] _RAND_850;
  reg [31:0] _RAND_851;
  reg [31:0] _RAND_852;
  reg [31:0] _RAND_853;
  reg [31:0] _RAND_854;
  reg [31:0] _RAND_855;
  reg [31:0] _RAND_856;
  reg [31:0] _RAND_857;
  reg [31:0] _RAND_858;
  reg [31:0] _RAND_859;
  reg [31:0] _RAND_860;
  reg [31:0] _RAND_861;
  reg [31:0] _RAND_862;
  reg [31:0] _RAND_863;
  reg [31:0] _RAND_864;
  reg [31:0] _RAND_865;
  reg [31:0] _RAND_866;
  reg [31:0] _RAND_867;
  reg [31:0] _RAND_868;
  reg [31:0] _RAND_869;
  reg [31:0] _RAND_870;
  reg [31:0] _RAND_871;
  reg [31:0] _RAND_872;
  reg [31:0] _RAND_873;
  reg [31:0] _RAND_874;
  reg [31:0] _RAND_875;
  reg [31:0] _RAND_876;
  reg [31:0] _RAND_877;
  reg [31:0] _RAND_878;
  reg [31:0] _RAND_879;
  reg [31:0] _RAND_880;
  reg [31:0] _RAND_881;
  reg [31:0] _RAND_882;
  reg [31:0] _RAND_883;
  reg [31:0] _RAND_884;
  reg [31:0] _RAND_885;
  reg [31:0] _RAND_886;
  reg [31:0] _RAND_887;
  reg [31:0] _RAND_888;
  reg [31:0] _RAND_889;
  reg [31:0] _RAND_890;
  reg [31:0] _RAND_891;
  reg [31:0] _RAND_892;
  reg [31:0] _RAND_893;
  reg [31:0] _RAND_894;
  reg [31:0] _RAND_895;
  reg [31:0] _RAND_896;
  reg [31:0] _RAND_897;
`endif // RANDOMIZE_REG_INIT
  wire [127:0] req_Q; // @[DCache.scala 225:19]
  wire  req_CLK; // @[DCache.scala 225:19]
  wire  req_CEN; // @[DCache.scala 225:19]
  wire  req_WEN; // @[DCache.scala 225:19]
  wire [127:0] req_BWEN; // @[DCache.scala 225:19]
  wire [7:0] req_A; // @[DCache.scala 225:19]
  wire [127:0] req_D; // @[DCache.scala 225:19]
  reg  way0V_0; // @[DCache.scala 33:22]
  reg  way0V_1; // @[DCache.scala 33:22]
  reg  way0V_2; // @[DCache.scala 33:22]
  reg  way0V_3; // @[DCache.scala 33:22]
  reg  way0V_4; // @[DCache.scala 33:22]
  reg  way0V_5; // @[DCache.scala 33:22]
  reg  way0V_6; // @[DCache.scala 33:22]
  reg  way0V_7; // @[DCache.scala 33:22]
  reg  way0V_8; // @[DCache.scala 33:22]
  reg  way0V_9; // @[DCache.scala 33:22]
  reg  way0V_10; // @[DCache.scala 33:22]
  reg  way0V_11; // @[DCache.scala 33:22]
  reg  way0V_12; // @[DCache.scala 33:22]
  reg  way0V_13; // @[DCache.scala 33:22]
  reg  way0V_14; // @[DCache.scala 33:22]
  reg  way0V_15; // @[DCache.scala 33:22]
  reg  way0V_16; // @[DCache.scala 33:22]
  reg  way0V_17; // @[DCache.scala 33:22]
  reg  way0V_18; // @[DCache.scala 33:22]
  reg  way0V_19; // @[DCache.scala 33:22]
  reg  way0V_20; // @[DCache.scala 33:22]
  reg  way0V_21; // @[DCache.scala 33:22]
  reg  way0V_22; // @[DCache.scala 33:22]
  reg  way0V_23; // @[DCache.scala 33:22]
  reg  way0V_24; // @[DCache.scala 33:22]
  reg  way0V_25; // @[DCache.scala 33:22]
  reg  way0V_26; // @[DCache.scala 33:22]
  reg  way0V_27; // @[DCache.scala 33:22]
  reg  way0V_28; // @[DCache.scala 33:22]
  reg  way0V_29; // @[DCache.scala 33:22]
  reg  way0V_30; // @[DCache.scala 33:22]
  reg  way0V_31; // @[DCache.scala 33:22]
  reg  way0V_32; // @[DCache.scala 33:22]
  reg  way0V_33; // @[DCache.scala 33:22]
  reg  way0V_34; // @[DCache.scala 33:22]
  reg  way0V_35; // @[DCache.scala 33:22]
  reg  way0V_36; // @[DCache.scala 33:22]
  reg  way0V_37; // @[DCache.scala 33:22]
  reg  way0V_38; // @[DCache.scala 33:22]
  reg  way0V_39; // @[DCache.scala 33:22]
  reg  way0V_40; // @[DCache.scala 33:22]
  reg  way0V_41; // @[DCache.scala 33:22]
  reg  way0V_42; // @[DCache.scala 33:22]
  reg  way0V_43; // @[DCache.scala 33:22]
  reg  way0V_44; // @[DCache.scala 33:22]
  reg  way0V_45; // @[DCache.scala 33:22]
  reg  way0V_46; // @[DCache.scala 33:22]
  reg  way0V_47; // @[DCache.scala 33:22]
  reg  way0V_48; // @[DCache.scala 33:22]
  reg  way0V_49; // @[DCache.scala 33:22]
  reg  way0V_50; // @[DCache.scala 33:22]
  reg  way0V_51; // @[DCache.scala 33:22]
  reg  way0V_52; // @[DCache.scala 33:22]
  reg  way0V_53; // @[DCache.scala 33:22]
  reg  way0V_54; // @[DCache.scala 33:22]
  reg  way0V_55; // @[DCache.scala 33:22]
  reg  way0V_56; // @[DCache.scala 33:22]
  reg  way0V_57; // @[DCache.scala 33:22]
  reg  way0V_58; // @[DCache.scala 33:22]
  reg  way0V_59; // @[DCache.scala 33:22]
  reg  way0V_60; // @[DCache.scala 33:22]
  reg  way0V_61; // @[DCache.scala 33:22]
  reg  way0V_62; // @[DCache.scala 33:22]
  reg  way0V_63; // @[DCache.scala 33:22]
  reg  way0V_64; // @[DCache.scala 33:22]
  reg  way0V_65; // @[DCache.scala 33:22]
  reg  way0V_66; // @[DCache.scala 33:22]
  reg  way0V_67; // @[DCache.scala 33:22]
  reg  way0V_68; // @[DCache.scala 33:22]
  reg  way0V_69; // @[DCache.scala 33:22]
  reg  way0V_70; // @[DCache.scala 33:22]
  reg  way0V_71; // @[DCache.scala 33:22]
  reg  way0V_72; // @[DCache.scala 33:22]
  reg  way0V_73; // @[DCache.scala 33:22]
  reg  way0V_74; // @[DCache.scala 33:22]
  reg  way0V_75; // @[DCache.scala 33:22]
  reg  way0V_76; // @[DCache.scala 33:22]
  reg  way0V_77; // @[DCache.scala 33:22]
  reg  way0V_78; // @[DCache.scala 33:22]
  reg  way0V_79; // @[DCache.scala 33:22]
  reg  way0V_80; // @[DCache.scala 33:22]
  reg  way0V_81; // @[DCache.scala 33:22]
  reg  way0V_82; // @[DCache.scala 33:22]
  reg  way0V_83; // @[DCache.scala 33:22]
  reg  way0V_84; // @[DCache.scala 33:22]
  reg  way0V_85; // @[DCache.scala 33:22]
  reg  way0V_86; // @[DCache.scala 33:22]
  reg  way0V_87; // @[DCache.scala 33:22]
  reg  way0V_88; // @[DCache.scala 33:22]
  reg  way0V_89; // @[DCache.scala 33:22]
  reg  way0V_90; // @[DCache.scala 33:22]
  reg  way0V_91; // @[DCache.scala 33:22]
  reg  way0V_92; // @[DCache.scala 33:22]
  reg  way0V_93; // @[DCache.scala 33:22]
  reg  way0V_94; // @[DCache.scala 33:22]
  reg  way0V_95; // @[DCache.scala 33:22]
  reg  way0V_96; // @[DCache.scala 33:22]
  reg  way0V_97; // @[DCache.scala 33:22]
  reg  way0V_98; // @[DCache.scala 33:22]
  reg  way0V_99; // @[DCache.scala 33:22]
  reg  way0V_100; // @[DCache.scala 33:22]
  reg  way0V_101; // @[DCache.scala 33:22]
  reg  way0V_102; // @[DCache.scala 33:22]
  reg  way0V_103; // @[DCache.scala 33:22]
  reg  way0V_104; // @[DCache.scala 33:22]
  reg  way0V_105; // @[DCache.scala 33:22]
  reg  way0V_106; // @[DCache.scala 33:22]
  reg  way0V_107; // @[DCache.scala 33:22]
  reg  way0V_108; // @[DCache.scala 33:22]
  reg  way0V_109; // @[DCache.scala 33:22]
  reg  way0V_110; // @[DCache.scala 33:22]
  reg  way0V_111; // @[DCache.scala 33:22]
  reg  way0V_112; // @[DCache.scala 33:22]
  reg  way0V_113; // @[DCache.scala 33:22]
  reg  way0V_114; // @[DCache.scala 33:22]
  reg  way0V_115; // @[DCache.scala 33:22]
  reg  way0V_116; // @[DCache.scala 33:22]
  reg  way0V_117; // @[DCache.scala 33:22]
  reg  way0V_118; // @[DCache.scala 33:22]
  reg  way0V_119; // @[DCache.scala 33:22]
  reg  way0V_120; // @[DCache.scala 33:22]
  reg  way0V_121; // @[DCache.scala 33:22]
  reg  way0V_122; // @[DCache.scala 33:22]
  reg  way0V_123; // @[DCache.scala 33:22]
  reg  way0V_124; // @[DCache.scala 33:22]
  reg  way0V_125; // @[DCache.scala 33:22]
  reg  way0V_126; // @[DCache.scala 33:22]
  reg  way0V_127; // @[DCache.scala 33:22]
  reg [20:0] way0Tag_0; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_1; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_2; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_3; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_4; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_5; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_6; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_7; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_8; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_9; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_10; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_11; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_12; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_13; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_14; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_15; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_16; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_17; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_18; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_19; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_20; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_21; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_22; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_23; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_24; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_25; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_26; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_27; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_28; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_29; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_30; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_31; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_32; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_33; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_34; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_35; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_36; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_37; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_38; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_39; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_40; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_41; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_42; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_43; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_44; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_45; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_46; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_47; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_48; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_49; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_50; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_51; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_52; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_53; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_54; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_55; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_56; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_57; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_58; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_59; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_60; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_61; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_62; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_63; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_64; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_65; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_66; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_67; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_68; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_69; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_70; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_71; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_72; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_73; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_74; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_75; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_76; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_77; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_78; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_79; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_80; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_81; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_82; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_83; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_84; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_85; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_86; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_87; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_88; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_89; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_90; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_91; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_92; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_93; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_94; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_95; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_96; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_97; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_98; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_99; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_100; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_101; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_102; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_103; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_104; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_105; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_106; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_107; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_108; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_109; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_110; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_111; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_112; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_113; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_114; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_115; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_116; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_117; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_118; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_119; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_120; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_121; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_122; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_123; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_124; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_125; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_126; // @[DCache.scala 34:24]
  reg [20:0] way0Tag_127; // @[DCache.scala 34:24]
  reg  way0Age_0; // @[DCache.scala 36:24]
  reg  way0Age_1; // @[DCache.scala 36:24]
  reg  way0Age_2; // @[DCache.scala 36:24]
  reg  way0Age_3; // @[DCache.scala 36:24]
  reg  way0Age_4; // @[DCache.scala 36:24]
  reg  way0Age_5; // @[DCache.scala 36:24]
  reg  way0Age_6; // @[DCache.scala 36:24]
  reg  way0Age_7; // @[DCache.scala 36:24]
  reg  way0Age_8; // @[DCache.scala 36:24]
  reg  way0Age_9; // @[DCache.scala 36:24]
  reg  way0Age_10; // @[DCache.scala 36:24]
  reg  way0Age_11; // @[DCache.scala 36:24]
  reg  way0Age_12; // @[DCache.scala 36:24]
  reg  way0Age_13; // @[DCache.scala 36:24]
  reg  way0Age_14; // @[DCache.scala 36:24]
  reg  way0Age_15; // @[DCache.scala 36:24]
  reg  way0Age_16; // @[DCache.scala 36:24]
  reg  way0Age_17; // @[DCache.scala 36:24]
  reg  way0Age_18; // @[DCache.scala 36:24]
  reg  way0Age_19; // @[DCache.scala 36:24]
  reg  way0Age_20; // @[DCache.scala 36:24]
  reg  way0Age_21; // @[DCache.scala 36:24]
  reg  way0Age_22; // @[DCache.scala 36:24]
  reg  way0Age_23; // @[DCache.scala 36:24]
  reg  way0Age_24; // @[DCache.scala 36:24]
  reg  way0Age_25; // @[DCache.scala 36:24]
  reg  way0Age_26; // @[DCache.scala 36:24]
  reg  way0Age_27; // @[DCache.scala 36:24]
  reg  way0Age_28; // @[DCache.scala 36:24]
  reg  way0Age_29; // @[DCache.scala 36:24]
  reg  way0Age_30; // @[DCache.scala 36:24]
  reg  way0Age_31; // @[DCache.scala 36:24]
  reg  way0Age_32; // @[DCache.scala 36:24]
  reg  way0Age_33; // @[DCache.scala 36:24]
  reg  way0Age_34; // @[DCache.scala 36:24]
  reg  way0Age_35; // @[DCache.scala 36:24]
  reg  way0Age_36; // @[DCache.scala 36:24]
  reg  way0Age_37; // @[DCache.scala 36:24]
  reg  way0Age_38; // @[DCache.scala 36:24]
  reg  way0Age_39; // @[DCache.scala 36:24]
  reg  way0Age_40; // @[DCache.scala 36:24]
  reg  way0Age_41; // @[DCache.scala 36:24]
  reg  way0Age_42; // @[DCache.scala 36:24]
  reg  way0Age_43; // @[DCache.scala 36:24]
  reg  way0Age_44; // @[DCache.scala 36:24]
  reg  way0Age_45; // @[DCache.scala 36:24]
  reg  way0Age_46; // @[DCache.scala 36:24]
  reg  way0Age_47; // @[DCache.scala 36:24]
  reg  way0Age_48; // @[DCache.scala 36:24]
  reg  way0Age_49; // @[DCache.scala 36:24]
  reg  way0Age_50; // @[DCache.scala 36:24]
  reg  way0Age_51; // @[DCache.scala 36:24]
  reg  way0Age_52; // @[DCache.scala 36:24]
  reg  way0Age_53; // @[DCache.scala 36:24]
  reg  way0Age_54; // @[DCache.scala 36:24]
  reg  way0Age_55; // @[DCache.scala 36:24]
  reg  way0Age_56; // @[DCache.scala 36:24]
  reg  way0Age_57; // @[DCache.scala 36:24]
  reg  way0Age_58; // @[DCache.scala 36:24]
  reg  way0Age_59; // @[DCache.scala 36:24]
  reg  way0Age_60; // @[DCache.scala 36:24]
  reg  way0Age_61; // @[DCache.scala 36:24]
  reg  way0Age_62; // @[DCache.scala 36:24]
  reg  way0Age_63; // @[DCache.scala 36:24]
  reg  way0Age_64; // @[DCache.scala 36:24]
  reg  way0Age_65; // @[DCache.scala 36:24]
  reg  way0Age_66; // @[DCache.scala 36:24]
  reg  way0Age_67; // @[DCache.scala 36:24]
  reg  way0Age_68; // @[DCache.scala 36:24]
  reg  way0Age_69; // @[DCache.scala 36:24]
  reg  way0Age_70; // @[DCache.scala 36:24]
  reg  way0Age_71; // @[DCache.scala 36:24]
  reg  way0Age_72; // @[DCache.scala 36:24]
  reg  way0Age_73; // @[DCache.scala 36:24]
  reg  way0Age_74; // @[DCache.scala 36:24]
  reg  way0Age_75; // @[DCache.scala 36:24]
  reg  way0Age_76; // @[DCache.scala 36:24]
  reg  way0Age_77; // @[DCache.scala 36:24]
  reg  way0Age_78; // @[DCache.scala 36:24]
  reg  way0Age_79; // @[DCache.scala 36:24]
  reg  way0Age_80; // @[DCache.scala 36:24]
  reg  way0Age_81; // @[DCache.scala 36:24]
  reg  way0Age_82; // @[DCache.scala 36:24]
  reg  way0Age_83; // @[DCache.scala 36:24]
  reg  way0Age_84; // @[DCache.scala 36:24]
  reg  way0Age_85; // @[DCache.scala 36:24]
  reg  way0Age_86; // @[DCache.scala 36:24]
  reg  way0Age_87; // @[DCache.scala 36:24]
  reg  way0Age_88; // @[DCache.scala 36:24]
  reg  way0Age_89; // @[DCache.scala 36:24]
  reg  way0Age_90; // @[DCache.scala 36:24]
  reg  way0Age_91; // @[DCache.scala 36:24]
  reg  way0Age_92; // @[DCache.scala 36:24]
  reg  way0Age_93; // @[DCache.scala 36:24]
  reg  way0Age_94; // @[DCache.scala 36:24]
  reg  way0Age_95; // @[DCache.scala 36:24]
  reg  way0Age_96; // @[DCache.scala 36:24]
  reg  way0Age_97; // @[DCache.scala 36:24]
  reg  way0Age_98; // @[DCache.scala 36:24]
  reg  way0Age_99; // @[DCache.scala 36:24]
  reg  way0Age_100; // @[DCache.scala 36:24]
  reg  way0Age_101; // @[DCache.scala 36:24]
  reg  way0Age_102; // @[DCache.scala 36:24]
  reg  way0Age_103; // @[DCache.scala 36:24]
  reg  way0Age_104; // @[DCache.scala 36:24]
  reg  way0Age_105; // @[DCache.scala 36:24]
  reg  way0Age_106; // @[DCache.scala 36:24]
  reg  way0Age_107; // @[DCache.scala 36:24]
  reg  way0Age_108; // @[DCache.scala 36:24]
  reg  way0Age_109; // @[DCache.scala 36:24]
  reg  way0Age_110; // @[DCache.scala 36:24]
  reg  way0Age_111; // @[DCache.scala 36:24]
  reg  way0Age_112; // @[DCache.scala 36:24]
  reg  way0Age_113; // @[DCache.scala 36:24]
  reg  way0Age_114; // @[DCache.scala 36:24]
  reg  way0Age_115; // @[DCache.scala 36:24]
  reg  way0Age_116; // @[DCache.scala 36:24]
  reg  way0Age_117; // @[DCache.scala 36:24]
  reg  way0Age_118; // @[DCache.scala 36:24]
  reg  way0Age_119; // @[DCache.scala 36:24]
  reg  way0Age_120; // @[DCache.scala 36:24]
  reg  way0Age_121; // @[DCache.scala 36:24]
  reg  way0Age_122; // @[DCache.scala 36:24]
  reg  way0Age_123; // @[DCache.scala 36:24]
  reg  way0Age_124; // @[DCache.scala 36:24]
  reg  way0Age_125; // @[DCache.scala 36:24]
  reg  way0Age_126; // @[DCache.scala 36:24]
  reg  way0Age_127; // @[DCache.scala 36:24]
  reg  way0Dirty_0; // @[DCache.scala 37:26]
  reg  way0Dirty_1; // @[DCache.scala 37:26]
  reg  way0Dirty_2; // @[DCache.scala 37:26]
  reg  way0Dirty_3; // @[DCache.scala 37:26]
  reg  way0Dirty_4; // @[DCache.scala 37:26]
  reg  way0Dirty_5; // @[DCache.scala 37:26]
  reg  way0Dirty_6; // @[DCache.scala 37:26]
  reg  way0Dirty_7; // @[DCache.scala 37:26]
  reg  way0Dirty_8; // @[DCache.scala 37:26]
  reg  way0Dirty_9; // @[DCache.scala 37:26]
  reg  way0Dirty_10; // @[DCache.scala 37:26]
  reg  way0Dirty_11; // @[DCache.scala 37:26]
  reg  way0Dirty_12; // @[DCache.scala 37:26]
  reg  way0Dirty_13; // @[DCache.scala 37:26]
  reg  way0Dirty_14; // @[DCache.scala 37:26]
  reg  way0Dirty_15; // @[DCache.scala 37:26]
  reg  way0Dirty_16; // @[DCache.scala 37:26]
  reg  way0Dirty_17; // @[DCache.scala 37:26]
  reg  way0Dirty_18; // @[DCache.scala 37:26]
  reg  way0Dirty_19; // @[DCache.scala 37:26]
  reg  way0Dirty_20; // @[DCache.scala 37:26]
  reg  way0Dirty_21; // @[DCache.scala 37:26]
  reg  way0Dirty_22; // @[DCache.scala 37:26]
  reg  way0Dirty_23; // @[DCache.scala 37:26]
  reg  way0Dirty_24; // @[DCache.scala 37:26]
  reg  way0Dirty_25; // @[DCache.scala 37:26]
  reg  way0Dirty_26; // @[DCache.scala 37:26]
  reg  way0Dirty_27; // @[DCache.scala 37:26]
  reg  way0Dirty_28; // @[DCache.scala 37:26]
  reg  way0Dirty_29; // @[DCache.scala 37:26]
  reg  way0Dirty_30; // @[DCache.scala 37:26]
  reg  way0Dirty_31; // @[DCache.scala 37:26]
  reg  way0Dirty_32; // @[DCache.scala 37:26]
  reg  way0Dirty_33; // @[DCache.scala 37:26]
  reg  way0Dirty_34; // @[DCache.scala 37:26]
  reg  way0Dirty_35; // @[DCache.scala 37:26]
  reg  way0Dirty_36; // @[DCache.scala 37:26]
  reg  way0Dirty_37; // @[DCache.scala 37:26]
  reg  way0Dirty_38; // @[DCache.scala 37:26]
  reg  way0Dirty_39; // @[DCache.scala 37:26]
  reg  way0Dirty_40; // @[DCache.scala 37:26]
  reg  way0Dirty_41; // @[DCache.scala 37:26]
  reg  way0Dirty_42; // @[DCache.scala 37:26]
  reg  way0Dirty_43; // @[DCache.scala 37:26]
  reg  way0Dirty_44; // @[DCache.scala 37:26]
  reg  way0Dirty_45; // @[DCache.scala 37:26]
  reg  way0Dirty_46; // @[DCache.scala 37:26]
  reg  way0Dirty_47; // @[DCache.scala 37:26]
  reg  way0Dirty_48; // @[DCache.scala 37:26]
  reg  way0Dirty_49; // @[DCache.scala 37:26]
  reg  way0Dirty_50; // @[DCache.scala 37:26]
  reg  way0Dirty_51; // @[DCache.scala 37:26]
  reg  way0Dirty_52; // @[DCache.scala 37:26]
  reg  way0Dirty_53; // @[DCache.scala 37:26]
  reg  way0Dirty_54; // @[DCache.scala 37:26]
  reg  way0Dirty_55; // @[DCache.scala 37:26]
  reg  way0Dirty_56; // @[DCache.scala 37:26]
  reg  way0Dirty_57; // @[DCache.scala 37:26]
  reg  way0Dirty_58; // @[DCache.scala 37:26]
  reg  way0Dirty_59; // @[DCache.scala 37:26]
  reg  way0Dirty_60; // @[DCache.scala 37:26]
  reg  way0Dirty_61; // @[DCache.scala 37:26]
  reg  way0Dirty_62; // @[DCache.scala 37:26]
  reg  way0Dirty_63; // @[DCache.scala 37:26]
  reg  way0Dirty_64; // @[DCache.scala 37:26]
  reg  way0Dirty_65; // @[DCache.scala 37:26]
  reg  way0Dirty_66; // @[DCache.scala 37:26]
  reg  way0Dirty_67; // @[DCache.scala 37:26]
  reg  way0Dirty_68; // @[DCache.scala 37:26]
  reg  way0Dirty_69; // @[DCache.scala 37:26]
  reg  way0Dirty_70; // @[DCache.scala 37:26]
  reg  way0Dirty_71; // @[DCache.scala 37:26]
  reg  way0Dirty_72; // @[DCache.scala 37:26]
  reg  way0Dirty_73; // @[DCache.scala 37:26]
  reg  way0Dirty_74; // @[DCache.scala 37:26]
  reg  way0Dirty_75; // @[DCache.scala 37:26]
  reg  way0Dirty_76; // @[DCache.scala 37:26]
  reg  way0Dirty_77; // @[DCache.scala 37:26]
  reg  way0Dirty_78; // @[DCache.scala 37:26]
  reg  way0Dirty_79; // @[DCache.scala 37:26]
  reg  way0Dirty_80; // @[DCache.scala 37:26]
  reg  way0Dirty_81; // @[DCache.scala 37:26]
  reg  way0Dirty_82; // @[DCache.scala 37:26]
  reg  way0Dirty_83; // @[DCache.scala 37:26]
  reg  way0Dirty_84; // @[DCache.scala 37:26]
  reg  way0Dirty_85; // @[DCache.scala 37:26]
  reg  way0Dirty_86; // @[DCache.scala 37:26]
  reg  way0Dirty_87; // @[DCache.scala 37:26]
  reg  way0Dirty_88; // @[DCache.scala 37:26]
  reg  way0Dirty_89; // @[DCache.scala 37:26]
  reg  way0Dirty_90; // @[DCache.scala 37:26]
  reg  way0Dirty_91; // @[DCache.scala 37:26]
  reg  way0Dirty_92; // @[DCache.scala 37:26]
  reg  way0Dirty_93; // @[DCache.scala 37:26]
  reg  way0Dirty_94; // @[DCache.scala 37:26]
  reg  way0Dirty_95; // @[DCache.scala 37:26]
  reg  way0Dirty_96; // @[DCache.scala 37:26]
  reg  way0Dirty_97; // @[DCache.scala 37:26]
  reg  way0Dirty_98; // @[DCache.scala 37:26]
  reg  way0Dirty_99; // @[DCache.scala 37:26]
  reg  way0Dirty_100; // @[DCache.scala 37:26]
  reg  way0Dirty_101; // @[DCache.scala 37:26]
  reg  way0Dirty_102; // @[DCache.scala 37:26]
  reg  way0Dirty_103; // @[DCache.scala 37:26]
  reg  way0Dirty_104; // @[DCache.scala 37:26]
  reg  way0Dirty_105; // @[DCache.scala 37:26]
  reg  way0Dirty_106; // @[DCache.scala 37:26]
  reg  way0Dirty_107; // @[DCache.scala 37:26]
  reg  way0Dirty_108; // @[DCache.scala 37:26]
  reg  way0Dirty_109; // @[DCache.scala 37:26]
  reg  way0Dirty_110; // @[DCache.scala 37:26]
  reg  way0Dirty_111; // @[DCache.scala 37:26]
  reg  way0Dirty_112; // @[DCache.scala 37:26]
  reg  way0Dirty_113; // @[DCache.scala 37:26]
  reg  way0Dirty_114; // @[DCache.scala 37:26]
  reg  way0Dirty_115; // @[DCache.scala 37:26]
  reg  way0Dirty_116; // @[DCache.scala 37:26]
  reg  way0Dirty_117; // @[DCache.scala 37:26]
  reg  way0Dirty_118; // @[DCache.scala 37:26]
  reg  way0Dirty_119; // @[DCache.scala 37:26]
  reg  way0Dirty_120; // @[DCache.scala 37:26]
  reg  way0Dirty_121; // @[DCache.scala 37:26]
  reg  way0Dirty_122; // @[DCache.scala 37:26]
  reg  way0Dirty_123; // @[DCache.scala 37:26]
  reg  way0Dirty_124; // @[DCache.scala 37:26]
  reg  way0Dirty_125; // @[DCache.scala 37:26]
  reg  way0Dirty_126; // @[DCache.scala 37:26]
  reg  way0Dirty_127; // @[DCache.scala 37:26]
  reg  way1V_0; // @[DCache.scala 39:22]
  reg  way1V_1; // @[DCache.scala 39:22]
  reg  way1V_2; // @[DCache.scala 39:22]
  reg  way1V_3; // @[DCache.scala 39:22]
  reg  way1V_4; // @[DCache.scala 39:22]
  reg  way1V_5; // @[DCache.scala 39:22]
  reg  way1V_6; // @[DCache.scala 39:22]
  reg  way1V_7; // @[DCache.scala 39:22]
  reg  way1V_8; // @[DCache.scala 39:22]
  reg  way1V_9; // @[DCache.scala 39:22]
  reg  way1V_10; // @[DCache.scala 39:22]
  reg  way1V_11; // @[DCache.scala 39:22]
  reg  way1V_12; // @[DCache.scala 39:22]
  reg  way1V_13; // @[DCache.scala 39:22]
  reg  way1V_14; // @[DCache.scala 39:22]
  reg  way1V_15; // @[DCache.scala 39:22]
  reg  way1V_16; // @[DCache.scala 39:22]
  reg  way1V_17; // @[DCache.scala 39:22]
  reg  way1V_18; // @[DCache.scala 39:22]
  reg  way1V_19; // @[DCache.scala 39:22]
  reg  way1V_20; // @[DCache.scala 39:22]
  reg  way1V_21; // @[DCache.scala 39:22]
  reg  way1V_22; // @[DCache.scala 39:22]
  reg  way1V_23; // @[DCache.scala 39:22]
  reg  way1V_24; // @[DCache.scala 39:22]
  reg  way1V_25; // @[DCache.scala 39:22]
  reg  way1V_26; // @[DCache.scala 39:22]
  reg  way1V_27; // @[DCache.scala 39:22]
  reg  way1V_28; // @[DCache.scala 39:22]
  reg  way1V_29; // @[DCache.scala 39:22]
  reg  way1V_30; // @[DCache.scala 39:22]
  reg  way1V_31; // @[DCache.scala 39:22]
  reg  way1V_32; // @[DCache.scala 39:22]
  reg  way1V_33; // @[DCache.scala 39:22]
  reg  way1V_34; // @[DCache.scala 39:22]
  reg  way1V_35; // @[DCache.scala 39:22]
  reg  way1V_36; // @[DCache.scala 39:22]
  reg  way1V_37; // @[DCache.scala 39:22]
  reg  way1V_38; // @[DCache.scala 39:22]
  reg  way1V_39; // @[DCache.scala 39:22]
  reg  way1V_40; // @[DCache.scala 39:22]
  reg  way1V_41; // @[DCache.scala 39:22]
  reg  way1V_42; // @[DCache.scala 39:22]
  reg  way1V_43; // @[DCache.scala 39:22]
  reg  way1V_44; // @[DCache.scala 39:22]
  reg  way1V_45; // @[DCache.scala 39:22]
  reg  way1V_46; // @[DCache.scala 39:22]
  reg  way1V_47; // @[DCache.scala 39:22]
  reg  way1V_48; // @[DCache.scala 39:22]
  reg  way1V_49; // @[DCache.scala 39:22]
  reg  way1V_50; // @[DCache.scala 39:22]
  reg  way1V_51; // @[DCache.scala 39:22]
  reg  way1V_52; // @[DCache.scala 39:22]
  reg  way1V_53; // @[DCache.scala 39:22]
  reg  way1V_54; // @[DCache.scala 39:22]
  reg  way1V_55; // @[DCache.scala 39:22]
  reg  way1V_56; // @[DCache.scala 39:22]
  reg  way1V_57; // @[DCache.scala 39:22]
  reg  way1V_58; // @[DCache.scala 39:22]
  reg  way1V_59; // @[DCache.scala 39:22]
  reg  way1V_60; // @[DCache.scala 39:22]
  reg  way1V_61; // @[DCache.scala 39:22]
  reg  way1V_62; // @[DCache.scala 39:22]
  reg  way1V_63; // @[DCache.scala 39:22]
  reg  way1V_64; // @[DCache.scala 39:22]
  reg  way1V_65; // @[DCache.scala 39:22]
  reg  way1V_66; // @[DCache.scala 39:22]
  reg  way1V_67; // @[DCache.scala 39:22]
  reg  way1V_68; // @[DCache.scala 39:22]
  reg  way1V_69; // @[DCache.scala 39:22]
  reg  way1V_70; // @[DCache.scala 39:22]
  reg  way1V_71; // @[DCache.scala 39:22]
  reg  way1V_72; // @[DCache.scala 39:22]
  reg  way1V_73; // @[DCache.scala 39:22]
  reg  way1V_74; // @[DCache.scala 39:22]
  reg  way1V_75; // @[DCache.scala 39:22]
  reg  way1V_76; // @[DCache.scala 39:22]
  reg  way1V_77; // @[DCache.scala 39:22]
  reg  way1V_78; // @[DCache.scala 39:22]
  reg  way1V_79; // @[DCache.scala 39:22]
  reg  way1V_80; // @[DCache.scala 39:22]
  reg  way1V_81; // @[DCache.scala 39:22]
  reg  way1V_82; // @[DCache.scala 39:22]
  reg  way1V_83; // @[DCache.scala 39:22]
  reg  way1V_84; // @[DCache.scala 39:22]
  reg  way1V_85; // @[DCache.scala 39:22]
  reg  way1V_86; // @[DCache.scala 39:22]
  reg  way1V_87; // @[DCache.scala 39:22]
  reg  way1V_88; // @[DCache.scala 39:22]
  reg  way1V_89; // @[DCache.scala 39:22]
  reg  way1V_90; // @[DCache.scala 39:22]
  reg  way1V_91; // @[DCache.scala 39:22]
  reg  way1V_92; // @[DCache.scala 39:22]
  reg  way1V_93; // @[DCache.scala 39:22]
  reg  way1V_94; // @[DCache.scala 39:22]
  reg  way1V_95; // @[DCache.scala 39:22]
  reg  way1V_96; // @[DCache.scala 39:22]
  reg  way1V_97; // @[DCache.scala 39:22]
  reg  way1V_98; // @[DCache.scala 39:22]
  reg  way1V_99; // @[DCache.scala 39:22]
  reg  way1V_100; // @[DCache.scala 39:22]
  reg  way1V_101; // @[DCache.scala 39:22]
  reg  way1V_102; // @[DCache.scala 39:22]
  reg  way1V_103; // @[DCache.scala 39:22]
  reg  way1V_104; // @[DCache.scala 39:22]
  reg  way1V_105; // @[DCache.scala 39:22]
  reg  way1V_106; // @[DCache.scala 39:22]
  reg  way1V_107; // @[DCache.scala 39:22]
  reg  way1V_108; // @[DCache.scala 39:22]
  reg  way1V_109; // @[DCache.scala 39:22]
  reg  way1V_110; // @[DCache.scala 39:22]
  reg  way1V_111; // @[DCache.scala 39:22]
  reg  way1V_112; // @[DCache.scala 39:22]
  reg  way1V_113; // @[DCache.scala 39:22]
  reg  way1V_114; // @[DCache.scala 39:22]
  reg  way1V_115; // @[DCache.scala 39:22]
  reg  way1V_116; // @[DCache.scala 39:22]
  reg  way1V_117; // @[DCache.scala 39:22]
  reg  way1V_118; // @[DCache.scala 39:22]
  reg  way1V_119; // @[DCache.scala 39:22]
  reg  way1V_120; // @[DCache.scala 39:22]
  reg  way1V_121; // @[DCache.scala 39:22]
  reg  way1V_122; // @[DCache.scala 39:22]
  reg  way1V_123; // @[DCache.scala 39:22]
  reg  way1V_124; // @[DCache.scala 39:22]
  reg  way1V_125; // @[DCache.scala 39:22]
  reg  way1V_126; // @[DCache.scala 39:22]
  reg  way1V_127; // @[DCache.scala 39:22]
  reg [20:0] way1Tag_0; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_1; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_2; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_3; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_4; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_5; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_6; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_7; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_8; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_9; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_10; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_11; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_12; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_13; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_14; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_15; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_16; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_17; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_18; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_19; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_20; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_21; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_22; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_23; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_24; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_25; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_26; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_27; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_28; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_29; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_30; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_31; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_32; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_33; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_34; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_35; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_36; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_37; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_38; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_39; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_40; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_41; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_42; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_43; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_44; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_45; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_46; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_47; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_48; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_49; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_50; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_51; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_52; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_53; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_54; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_55; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_56; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_57; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_58; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_59; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_60; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_61; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_62; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_63; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_64; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_65; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_66; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_67; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_68; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_69; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_70; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_71; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_72; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_73; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_74; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_75; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_76; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_77; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_78; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_79; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_80; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_81; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_82; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_83; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_84; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_85; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_86; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_87; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_88; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_89; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_90; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_91; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_92; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_93; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_94; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_95; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_96; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_97; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_98; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_99; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_100; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_101; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_102; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_103; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_104; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_105; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_106; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_107; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_108; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_109; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_110; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_111; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_112; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_113; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_114; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_115; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_116; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_117; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_118; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_119; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_120; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_121; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_122; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_123; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_124; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_125; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_126; // @[DCache.scala 40:24]
  reg [20:0] way1Tag_127; // @[DCache.scala 40:24]
  reg  way1Dirty_0; // @[DCache.scala 43:26]
  reg  way1Dirty_1; // @[DCache.scala 43:26]
  reg  way1Dirty_2; // @[DCache.scala 43:26]
  reg  way1Dirty_3; // @[DCache.scala 43:26]
  reg  way1Dirty_4; // @[DCache.scala 43:26]
  reg  way1Dirty_5; // @[DCache.scala 43:26]
  reg  way1Dirty_6; // @[DCache.scala 43:26]
  reg  way1Dirty_7; // @[DCache.scala 43:26]
  reg  way1Dirty_8; // @[DCache.scala 43:26]
  reg  way1Dirty_9; // @[DCache.scala 43:26]
  reg  way1Dirty_10; // @[DCache.scala 43:26]
  reg  way1Dirty_11; // @[DCache.scala 43:26]
  reg  way1Dirty_12; // @[DCache.scala 43:26]
  reg  way1Dirty_13; // @[DCache.scala 43:26]
  reg  way1Dirty_14; // @[DCache.scala 43:26]
  reg  way1Dirty_15; // @[DCache.scala 43:26]
  reg  way1Dirty_16; // @[DCache.scala 43:26]
  reg  way1Dirty_17; // @[DCache.scala 43:26]
  reg  way1Dirty_18; // @[DCache.scala 43:26]
  reg  way1Dirty_19; // @[DCache.scala 43:26]
  reg  way1Dirty_20; // @[DCache.scala 43:26]
  reg  way1Dirty_21; // @[DCache.scala 43:26]
  reg  way1Dirty_22; // @[DCache.scala 43:26]
  reg  way1Dirty_23; // @[DCache.scala 43:26]
  reg  way1Dirty_24; // @[DCache.scala 43:26]
  reg  way1Dirty_25; // @[DCache.scala 43:26]
  reg  way1Dirty_26; // @[DCache.scala 43:26]
  reg  way1Dirty_27; // @[DCache.scala 43:26]
  reg  way1Dirty_28; // @[DCache.scala 43:26]
  reg  way1Dirty_29; // @[DCache.scala 43:26]
  reg  way1Dirty_30; // @[DCache.scala 43:26]
  reg  way1Dirty_31; // @[DCache.scala 43:26]
  reg  way1Dirty_32; // @[DCache.scala 43:26]
  reg  way1Dirty_33; // @[DCache.scala 43:26]
  reg  way1Dirty_34; // @[DCache.scala 43:26]
  reg  way1Dirty_35; // @[DCache.scala 43:26]
  reg  way1Dirty_36; // @[DCache.scala 43:26]
  reg  way1Dirty_37; // @[DCache.scala 43:26]
  reg  way1Dirty_38; // @[DCache.scala 43:26]
  reg  way1Dirty_39; // @[DCache.scala 43:26]
  reg  way1Dirty_40; // @[DCache.scala 43:26]
  reg  way1Dirty_41; // @[DCache.scala 43:26]
  reg  way1Dirty_42; // @[DCache.scala 43:26]
  reg  way1Dirty_43; // @[DCache.scala 43:26]
  reg  way1Dirty_44; // @[DCache.scala 43:26]
  reg  way1Dirty_45; // @[DCache.scala 43:26]
  reg  way1Dirty_46; // @[DCache.scala 43:26]
  reg  way1Dirty_47; // @[DCache.scala 43:26]
  reg  way1Dirty_48; // @[DCache.scala 43:26]
  reg  way1Dirty_49; // @[DCache.scala 43:26]
  reg  way1Dirty_50; // @[DCache.scala 43:26]
  reg  way1Dirty_51; // @[DCache.scala 43:26]
  reg  way1Dirty_52; // @[DCache.scala 43:26]
  reg  way1Dirty_53; // @[DCache.scala 43:26]
  reg  way1Dirty_54; // @[DCache.scala 43:26]
  reg  way1Dirty_55; // @[DCache.scala 43:26]
  reg  way1Dirty_56; // @[DCache.scala 43:26]
  reg  way1Dirty_57; // @[DCache.scala 43:26]
  reg  way1Dirty_58; // @[DCache.scala 43:26]
  reg  way1Dirty_59; // @[DCache.scala 43:26]
  reg  way1Dirty_60; // @[DCache.scala 43:26]
  reg  way1Dirty_61; // @[DCache.scala 43:26]
  reg  way1Dirty_62; // @[DCache.scala 43:26]
  reg  way1Dirty_63; // @[DCache.scala 43:26]
  reg  way1Dirty_64; // @[DCache.scala 43:26]
  reg  way1Dirty_65; // @[DCache.scala 43:26]
  reg  way1Dirty_66; // @[DCache.scala 43:26]
  reg  way1Dirty_67; // @[DCache.scala 43:26]
  reg  way1Dirty_68; // @[DCache.scala 43:26]
  reg  way1Dirty_69; // @[DCache.scala 43:26]
  reg  way1Dirty_70; // @[DCache.scala 43:26]
  reg  way1Dirty_71; // @[DCache.scala 43:26]
  reg  way1Dirty_72; // @[DCache.scala 43:26]
  reg  way1Dirty_73; // @[DCache.scala 43:26]
  reg  way1Dirty_74; // @[DCache.scala 43:26]
  reg  way1Dirty_75; // @[DCache.scala 43:26]
  reg  way1Dirty_76; // @[DCache.scala 43:26]
  reg  way1Dirty_77; // @[DCache.scala 43:26]
  reg  way1Dirty_78; // @[DCache.scala 43:26]
  reg  way1Dirty_79; // @[DCache.scala 43:26]
  reg  way1Dirty_80; // @[DCache.scala 43:26]
  reg  way1Dirty_81; // @[DCache.scala 43:26]
  reg  way1Dirty_82; // @[DCache.scala 43:26]
  reg  way1Dirty_83; // @[DCache.scala 43:26]
  reg  way1Dirty_84; // @[DCache.scala 43:26]
  reg  way1Dirty_85; // @[DCache.scala 43:26]
  reg  way1Dirty_86; // @[DCache.scala 43:26]
  reg  way1Dirty_87; // @[DCache.scala 43:26]
  reg  way1Dirty_88; // @[DCache.scala 43:26]
  reg  way1Dirty_89; // @[DCache.scala 43:26]
  reg  way1Dirty_90; // @[DCache.scala 43:26]
  reg  way1Dirty_91; // @[DCache.scala 43:26]
  reg  way1Dirty_92; // @[DCache.scala 43:26]
  reg  way1Dirty_93; // @[DCache.scala 43:26]
  reg  way1Dirty_94; // @[DCache.scala 43:26]
  reg  way1Dirty_95; // @[DCache.scala 43:26]
  reg  way1Dirty_96; // @[DCache.scala 43:26]
  reg  way1Dirty_97; // @[DCache.scala 43:26]
  reg  way1Dirty_98; // @[DCache.scala 43:26]
  reg  way1Dirty_99; // @[DCache.scala 43:26]
  reg  way1Dirty_100; // @[DCache.scala 43:26]
  reg  way1Dirty_101; // @[DCache.scala 43:26]
  reg  way1Dirty_102; // @[DCache.scala 43:26]
  reg  way1Dirty_103; // @[DCache.scala 43:26]
  reg  way1Dirty_104; // @[DCache.scala 43:26]
  reg  way1Dirty_105; // @[DCache.scala 43:26]
  reg  way1Dirty_106; // @[DCache.scala 43:26]
  reg  way1Dirty_107; // @[DCache.scala 43:26]
  reg  way1Dirty_108; // @[DCache.scala 43:26]
  reg  way1Dirty_109; // @[DCache.scala 43:26]
  reg  way1Dirty_110; // @[DCache.scala 43:26]
  reg  way1Dirty_111; // @[DCache.scala 43:26]
  reg  way1Dirty_112; // @[DCache.scala 43:26]
  reg  way1Dirty_113; // @[DCache.scala 43:26]
  reg  way1Dirty_114; // @[DCache.scala 43:26]
  reg  way1Dirty_115; // @[DCache.scala 43:26]
  reg  way1Dirty_116; // @[DCache.scala 43:26]
  reg  way1Dirty_117; // @[DCache.scala 43:26]
  reg  way1Dirty_118; // @[DCache.scala 43:26]
  reg  way1Dirty_119; // @[DCache.scala 43:26]
  reg  way1Dirty_120; // @[DCache.scala 43:26]
  reg  way1Dirty_121; // @[DCache.scala 43:26]
  reg  way1Dirty_122; // @[DCache.scala 43:26]
  reg  way1Dirty_123; // @[DCache.scala 43:26]
  reg  way1Dirty_124; // @[DCache.scala 43:26]
  reg  way1Dirty_125; // @[DCache.scala 43:26]
  reg  way1Dirty_126; // @[DCache.scala 43:26]
  reg  way1Dirty_127; // @[DCache.scala 43:26]
  reg [2:0] state; // @[DCache.scala 46:22]
  wire [20:0] reqTag = io_dmem_data_addr[31:11]; // @[DCache.scala 50:25]
  wire [6:0] reqIndex = io_dmem_data_addr[10:4]; // @[DCache.scala 51:27]
  wire [3:0] reqOff = io_dmem_data_addr[3:0]; // @[DCache.scala 52:25]
  wire [7:0] _strbT_T_1 = 8'h1 == io_dmem_data_strb ? 8'hff : 8'h0; // @[Mux.scala 81:58]
  wire [15:0] _strbT_T_3 = 8'h2 == io_dmem_data_strb ? 16'hff00 : {{8'd0}, _strbT_T_1}; // @[Mux.scala 81:58]
  wire [23:0] _strbT_T_5 = 8'h4 == io_dmem_data_strb ? 24'hff0000 : {{8'd0}, _strbT_T_3}; // @[Mux.scala 81:58]
  wire [31:0] _strbT_T_7 = 8'h8 == io_dmem_data_strb ? 32'hff000000 : {{8'd0}, _strbT_T_5}; // @[Mux.scala 81:58]
  wire [39:0] _strbT_T_9 = 8'h10 == io_dmem_data_strb ? 40'hff00000000 : {{8'd0}, _strbT_T_7}; // @[Mux.scala 81:58]
  wire [47:0] _strbT_T_11 = 8'h20 == io_dmem_data_strb ? 48'hff0000000000 : {{8'd0}, _strbT_T_9}; // @[Mux.scala 81:58]
  wire [55:0] _strbT_T_13 = 8'h40 == io_dmem_data_strb ? 56'hff000000000000 : {{8'd0}, _strbT_T_11}; // @[Mux.scala 81:58]
  wire [63:0] _strbT_T_15 = 8'h80 == io_dmem_data_strb ? 64'hff00000000000000 : {{8'd0}, _strbT_T_13}; // @[Mux.scala 81:58]
  wire [63:0] _strbT_T_17 = 8'h3 == io_dmem_data_strb ? 64'hffff : _strbT_T_15; // @[Mux.scala 81:58]
  wire [63:0] _strbT_T_19 = 8'hc == io_dmem_data_strb ? 64'hffff0000 : _strbT_T_17; // @[Mux.scala 81:58]
  wire [63:0] _strbT_T_21 = 8'h30 == io_dmem_data_strb ? 64'hffff00000000 : _strbT_T_19; // @[Mux.scala 81:58]
  wire [63:0] _strbT_T_23 = 8'hc0 == io_dmem_data_strb ? 64'hffff000000000000 : _strbT_T_21; // @[Mux.scala 81:58]
  wire [63:0] _strbT_T_25 = 8'hf == io_dmem_data_strb ? 64'hffffffff : _strbT_T_23; // @[Mux.scala 81:58]
  wire [63:0] _strbT_T_27 = 8'hf0 == io_dmem_data_strb ? 64'hffffffff00000000 : _strbT_T_25; // @[Mux.scala 81:58]
  wire [63:0] strbT = 8'hff == io_dmem_data_strb ? 64'hffffffffffffffff : _strbT_T_27; // @[Mux.scala 81:58]
  wire [64:0] _valid_strb_T_1 = {strbT,1'h0}; // @[Cat.scala 31:58]
  wire [64:0] _valid_strb_T_2 = {1'h0,strbT}; // @[Cat.scala 31:58]
  wire [64:0] valid_strb = reqOff[3] ? _valid_strb_T_1 : _valid_strb_T_2; // @[DCache.scala 75:23]
  wire  _GEN_140 = 7'h1 == reqIndex ? way0V_1 : way0V_0; // @[DCache.scala 120:{33,33}]
  wire  _GEN_141 = 7'h2 == reqIndex ? way0V_2 : _GEN_140; // @[DCache.scala 120:{33,33}]
  wire  _GEN_142 = 7'h3 == reqIndex ? way0V_3 : _GEN_141; // @[DCache.scala 120:{33,33}]
  wire  _GEN_143 = 7'h4 == reqIndex ? way0V_4 : _GEN_142; // @[DCache.scala 120:{33,33}]
  wire  _GEN_144 = 7'h5 == reqIndex ? way0V_5 : _GEN_143; // @[DCache.scala 120:{33,33}]
  wire  _GEN_145 = 7'h6 == reqIndex ? way0V_6 : _GEN_144; // @[DCache.scala 120:{33,33}]
  wire  _GEN_146 = 7'h7 == reqIndex ? way0V_7 : _GEN_145; // @[DCache.scala 120:{33,33}]
  wire  _GEN_147 = 7'h8 == reqIndex ? way0V_8 : _GEN_146; // @[DCache.scala 120:{33,33}]
  wire  _GEN_148 = 7'h9 == reqIndex ? way0V_9 : _GEN_147; // @[DCache.scala 120:{33,33}]
  wire  _GEN_149 = 7'ha == reqIndex ? way0V_10 : _GEN_148; // @[DCache.scala 120:{33,33}]
  wire  _GEN_150 = 7'hb == reqIndex ? way0V_11 : _GEN_149; // @[DCache.scala 120:{33,33}]
  wire  _GEN_151 = 7'hc == reqIndex ? way0V_12 : _GEN_150; // @[DCache.scala 120:{33,33}]
  wire  _GEN_152 = 7'hd == reqIndex ? way0V_13 : _GEN_151; // @[DCache.scala 120:{33,33}]
  wire  _GEN_153 = 7'he == reqIndex ? way0V_14 : _GEN_152; // @[DCache.scala 120:{33,33}]
  wire  _GEN_154 = 7'hf == reqIndex ? way0V_15 : _GEN_153; // @[DCache.scala 120:{33,33}]
  wire  _GEN_155 = 7'h10 == reqIndex ? way0V_16 : _GEN_154; // @[DCache.scala 120:{33,33}]
  wire  _GEN_156 = 7'h11 == reqIndex ? way0V_17 : _GEN_155; // @[DCache.scala 120:{33,33}]
  wire  _GEN_157 = 7'h12 == reqIndex ? way0V_18 : _GEN_156; // @[DCache.scala 120:{33,33}]
  wire  _GEN_158 = 7'h13 == reqIndex ? way0V_19 : _GEN_157; // @[DCache.scala 120:{33,33}]
  wire  _GEN_159 = 7'h14 == reqIndex ? way0V_20 : _GEN_158; // @[DCache.scala 120:{33,33}]
  wire  _GEN_160 = 7'h15 == reqIndex ? way0V_21 : _GEN_159; // @[DCache.scala 120:{33,33}]
  wire  _GEN_161 = 7'h16 == reqIndex ? way0V_22 : _GEN_160; // @[DCache.scala 120:{33,33}]
  wire  _GEN_162 = 7'h17 == reqIndex ? way0V_23 : _GEN_161; // @[DCache.scala 120:{33,33}]
  wire  _GEN_163 = 7'h18 == reqIndex ? way0V_24 : _GEN_162; // @[DCache.scala 120:{33,33}]
  wire  _GEN_164 = 7'h19 == reqIndex ? way0V_25 : _GEN_163; // @[DCache.scala 120:{33,33}]
  wire  _GEN_165 = 7'h1a == reqIndex ? way0V_26 : _GEN_164; // @[DCache.scala 120:{33,33}]
  wire  _GEN_166 = 7'h1b == reqIndex ? way0V_27 : _GEN_165; // @[DCache.scala 120:{33,33}]
  wire  _GEN_167 = 7'h1c == reqIndex ? way0V_28 : _GEN_166; // @[DCache.scala 120:{33,33}]
  wire  _GEN_168 = 7'h1d == reqIndex ? way0V_29 : _GEN_167; // @[DCache.scala 120:{33,33}]
  wire  _GEN_169 = 7'h1e == reqIndex ? way0V_30 : _GEN_168; // @[DCache.scala 120:{33,33}]
  wire  _GEN_170 = 7'h1f == reqIndex ? way0V_31 : _GEN_169; // @[DCache.scala 120:{33,33}]
  wire  _GEN_171 = 7'h20 == reqIndex ? way0V_32 : _GEN_170; // @[DCache.scala 120:{33,33}]
  wire  _GEN_172 = 7'h21 == reqIndex ? way0V_33 : _GEN_171; // @[DCache.scala 120:{33,33}]
  wire  _GEN_173 = 7'h22 == reqIndex ? way0V_34 : _GEN_172; // @[DCache.scala 120:{33,33}]
  wire  _GEN_174 = 7'h23 == reqIndex ? way0V_35 : _GEN_173; // @[DCache.scala 120:{33,33}]
  wire  _GEN_175 = 7'h24 == reqIndex ? way0V_36 : _GEN_174; // @[DCache.scala 120:{33,33}]
  wire  _GEN_176 = 7'h25 == reqIndex ? way0V_37 : _GEN_175; // @[DCache.scala 120:{33,33}]
  wire  _GEN_177 = 7'h26 == reqIndex ? way0V_38 : _GEN_176; // @[DCache.scala 120:{33,33}]
  wire  _GEN_178 = 7'h27 == reqIndex ? way0V_39 : _GEN_177; // @[DCache.scala 120:{33,33}]
  wire  _GEN_179 = 7'h28 == reqIndex ? way0V_40 : _GEN_178; // @[DCache.scala 120:{33,33}]
  wire  _GEN_180 = 7'h29 == reqIndex ? way0V_41 : _GEN_179; // @[DCache.scala 120:{33,33}]
  wire  _GEN_181 = 7'h2a == reqIndex ? way0V_42 : _GEN_180; // @[DCache.scala 120:{33,33}]
  wire  _GEN_182 = 7'h2b == reqIndex ? way0V_43 : _GEN_181; // @[DCache.scala 120:{33,33}]
  wire  _GEN_183 = 7'h2c == reqIndex ? way0V_44 : _GEN_182; // @[DCache.scala 120:{33,33}]
  wire  _GEN_184 = 7'h2d == reqIndex ? way0V_45 : _GEN_183; // @[DCache.scala 120:{33,33}]
  wire  _GEN_185 = 7'h2e == reqIndex ? way0V_46 : _GEN_184; // @[DCache.scala 120:{33,33}]
  wire  _GEN_186 = 7'h2f == reqIndex ? way0V_47 : _GEN_185; // @[DCache.scala 120:{33,33}]
  wire  _GEN_187 = 7'h30 == reqIndex ? way0V_48 : _GEN_186; // @[DCache.scala 120:{33,33}]
  wire  _GEN_188 = 7'h31 == reqIndex ? way0V_49 : _GEN_187; // @[DCache.scala 120:{33,33}]
  wire  _GEN_189 = 7'h32 == reqIndex ? way0V_50 : _GEN_188; // @[DCache.scala 120:{33,33}]
  wire  _GEN_190 = 7'h33 == reqIndex ? way0V_51 : _GEN_189; // @[DCache.scala 120:{33,33}]
  wire  _GEN_191 = 7'h34 == reqIndex ? way0V_52 : _GEN_190; // @[DCache.scala 120:{33,33}]
  wire  _GEN_192 = 7'h35 == reqIndex ? way0V_53 : _GEN_191; // @[DCache.scala 120:{33,33}]
  wire  _GEN_193 = 7'h36 == reqIndex ? way0V_54 : _GEN_192; // @[DCache.scala 120:{33,33}]
  wire  _GEN_194 = 7'h37 == reqIndex ? way0V_55 : _GEN_193; // @[DCache.scala 120:{33,33}]
  wire  _GEN_195 = 7'h38 == reqIndex ? way0V_56 : _GEN_194; // @[DCache.scala 120:{33,33}]
  wire  _GEN_196 = 7'h39 == reqIndex ? way0V_57 : _GEN_195; // @[DCache.scala 120:{33,33}]
  wire  _GEN_197 = 7'h3a == reqIndex ? way0V_58 : _GEN_196; // @[DCache.scala 120:{33,33}]
  wire  _GEN_198 = 7'h3b == reqIndex ? way0V_59 : _GEN_197; // @[DCache.scala 120:{33,33}]
  wire  _GEN_199 = 7'h3c == reqIndex ? way0V_60 : _GEN_198; // @[DCache.scala 120:{33,33}]
  wire  _GEN_200 = 7'h3d == reqIndex ? way0V_61 : _GEN_199; // @[DCache.scala 120:{33,33}]
  wire  _GEN_201 = 7'h3e == reqIndex ? way0V_62 : _GEN_200; // @[DCache.scala 120:{33,33}]
  wire  _GEN_202 = 7'h3f == reqIndex ? way0V_63 : _GEN_201; // @[DCache.scala 120:{33,33}]
  wire  _GEN_203 = 7'h40 == reqIndex ? way0V_64 : _GEN_202; // @[DCache.scala 120:{33,33}]
  wire  _GEN_204 = 7'h41 == reqIndex ? way0V_65 : _GEN_203; // @[DCache.scala 120:{33,33}]
  wire  _GEN_205 = 7'h42 == reqIndex ? way0V_66 : _GEN_204; // @[DCache.scala 120:{33,33}]
  wire  _GEN_206 = 7'h43 == reqIndex ? way0V_67 : _GEN_205; // @[DCache.scala 120:{33,33}]
  wire  _GEN_207 = 7'h44 == reqIndex ? way0V_68 : _GEN_206; // @[DCache.scala 120:{33,33}]
  wire  _GEN_208 = 7'h45 == reqIndex ? way0V_69 : _GEN_207; // @[DCache.scala 120:{33,33}]
  wire  _GEN_209 = 7'h46 == reqIndex ? way0V_70 : _GEN_208; // @[DCache.scala 120:{33,33}]
  wire  _GEN_210 = 7'h47 == reqIndex ? way0V_71 : _GEN_209; // @[DCache.scala 120:{33,33}]
  wire  _GEN_211 = 7'h48 == reqIndex ? way0V_72 : _GEN_210; // @[DCache.scala 120:{33,33}]
  wire  _GEN_212 = 7'h49 == reqIndex ? way0V_73 : _GEN_211; // @[DCache.scala 120:{33,33}]
  wire  _GEN_213 = 7'h4a == reqIndex ? way0V_74 : _GEN_212; // @[DCache.scala 120:{33,33}]
  wire  _GEN_214 = 7'h4b == reqIndex ? way0V_75 : _GEN_213; // @[DCache.scala 120:{33,33}]
  wire  _GEN_215 = 7'h4c == reqIndex ? way0V_76 : _GEN_214; // @[DCache.scala 120:{33,33}]
  wire  _GEN_216 = 7'h4d == reqIndex ? way0V_77 : _GEN_215; // @[DCache.scala 120:{33,33}]
  wire  _GEN_217 = 7'h4e == reqIndex ? way0V_78 : _GEN_216; // @[DCache.scala 120:{33,33}]
  wire  _GEN_218 = 7'h4f == reqIndex ? way0V_79 : _GEN_217; // @[DCache.scala 120:{33,33}]
  wire  _GEN_219 = 7'h50 == reqIndex ? way0V_80 : _GEN_218; // @[DCache.scala 120:{33,33}]
  wire  _GEN_220 = 7'h51 == reqIndex ? way0V_81 : _GEN_219; // @[DCache.scala 120:{33,33}]
  wire  _GEN_221 = 7'h52 == reqIndex ? way0V_82 : _GEN_220; // @[DCache.scala 120:{33,33}]
  wire  _GEN_222 = 7'h53 == reqIndex ? way0V_83 : _GEN_221; // @[DCache.scala 120:{33,33}]
  wire  _GEN_223 = 7'h54 == reqIndex ? way0V_84 : _GEN_222; // @[DCache.scala 120:{33,33}]
  wire  _GEN_224 = 7'h55 == reqIndex ? way0V_85 : _GEN_223; // @[DCache.scala 120:{33,33}]
  wire  _GEN_225 = 7'h56 == reqIndex ? way0V_86 : _GEN_224; // @[DCache.scala 120:{33,33}]
  wire  _GEN_226 = 7'h57 == reqIndex ? way0V_87 : _GEN_225; // @[DCache.scala 120:{33,33}]
  wire  _GEN_227 = 7'h58 == reqIndex ? way0V_88 : _GEN_226; // @[DCache.scala 120:{33,33}]
  wire  _GEN_228 = 7'h59 == reqIndex ? way0V_89 : _GEN_227; // @[DCache.scala 120:{33,33}]
  wire  _GEN_229 = 7'h5a == reqIndex ? way0V_90 : _GEN_228; // @[DCache.scala 120:{33,33}]
  wire  _GEN_230 = 7'h5b == reqIndex ? way0V_91 : _GEN_229; // @[DCache.scala 120:{33,33}]
  wire  _GEN_231 = 7'h5c == reqIndex ? way0V_92 : _GEN_230; // @[DCache.scala 120:{33,33}]
  wire  _GEN_232 = 7'h5d == reqIndex ? way0V_93 : _GEN_231; // @[DCache.scala 120:{33,33}]
  wire  _GEN_233 = 7'h5e == reqIndex ? way0V_94 : _GEN_232; // @[DCache.scala 120:{33,33}]
  wire  _GEN_234 = 7'h5f == reqIndex ? way0V_95 : _GEN_233; // @[DCache.scala 120:{33,33}]
  wire  _GEN_235 = 7'h60 == reqIndex ? way0V_96 : _GEN_234; // @[DCache.scala 120:{33,33}]
  wire  _GEN_236 = 7'h61 == reqIndex ? way0V_97 : _GEN_235; // @[DCache.scala 120:{33,33}]
  wire  _GEN_237 = 7'h62 == reqIndex ? way0V_98 : _GEN_236; // @[DCache.scala 120:{33,33}]
  wire  _GEN_238 = 7'h63 == reqIndex ? way0V_99 : _GEN_237; // @[DCache.scala 120:{33,33}]
  wire  _GEN_239 = 7'h64 == reqIndex ? way0V_100 : _GEN_238; // @[DCache.scala 120:{33,33}]
  wire  _GEN_240 = 7'h65 == reqIndex ? way0V_101 : _GEN_239; // @[DCache.scala 120:{33,33}]
  wire  _GEN_241 = 7'h66 == reqIndex ? way0V_102 : _GEN_240; // @[DCache.scala 120:{33,33}]
  wire  _GEN_242 = 7'h67 == reqIndex ? way0V_103 : _GEN_241; // @[DCache.scala 120:{33,33}]
  wire  _GEN_243 = 7'h68 == reqIndex ? way0V_104 : _GEN_242; // @[DCache.scala 120:{33,33}]
  wire  _GEN_244 = 7'h69 == reqIndex ? way0V_105 : _GEN_243; // @[DCache.scala 120:{33,33}]
  wire  _GEN_245 = 7'h6a == reqIndex ? way0V_106 : _GEN_244; // @[DCache.scala 120:{33,33}]
  wire  _GEN_246 = 7'h6b == reqIndex ? way0V_107 : _GEN_245; // @[DCache.scala 120:{33,33}]
  wire  _GEN_247 = 7'h6c == reqIndex ? way0V_108 : _GEN_246; // @[DCache.scala 120:{33,33}]
  wire  _GEN_248 = 7'h6d == reqIndex ? way0V_109 : _GEN_247; // @[DCache.scala 120:{33,33}]
  wire  _GEN_249 = 7'h6e == reqIndex ? way0V_110 : _GEN_248; // @[DCache.scala 120:{33,33}]
  wire  _GEN_250 = 7'h6f == reqIndex ? way0V_111 : _GEN_249; // @[DCache.scala 120:{33,33}]
  wire  _GEN_251 = 7'h70 == reqIndex ? way0V_112 : _GEN_250; // @[DCache.scala 120:{33,33}]
  wire  _GEN_252 = 7'h71 == reqIndex ? way0V_113 : _GEN_251; // @[DCache.scala 120:{33,33}]
  wire  _GEN_253 = 7'h72 == reqIndex ? way0V_114 : _GEN_252; // @[DCache.scala 120:{33,33}]
  wire  _GEN_254 = 7'h73 == reqIndex ? way0V_115 : _GEN_253; // @[DCache.scala 120:{33,33}]
  wire  _GEN_255 = 7'h74 == reqIndex ? way0V_116 : _GEN_254; // @[DCache.scala 120:{33,33}]
  wire  _GEN_256 = 7'h75 == reqIndex ? way0V_117 : _GEN_255; // @[DCache.scala 120:{33,33}]
  wire  _GEN_257 = 7'h76 == reqIndex ? way0V_118 : _GEN_256; // @[DCache.scala 120:{33,33}]
  wire  _GEN_258 = 7'h77 == reqIndex ? way0V_119 : _GEN_257; // @[DCache.scala 120:{33,33}]
  wire  _GEN_259 = 7'h78 == reqIndex ? way0V_120 : _GEN_258; // @[DCache.scala 120:{33,33}]
  wire  _GEN_260 = 7'h79 == reqIndex ? way0V_121 : _GEN_259; // @[DCache.scala 120:{33,33}]
  wire  _GEN_261 = 7'h7a == reqIndex ? way0V_122 : _GEN_260; // @[DCache.scala 120:{33,33}]
  wire  _GEN_262 = 7'h7b == reqIndex ? way0V_123 : _GEN_261; // @[DCache.scala 120:{33,33}]
  wire  _GEN_263 = 7'h7c == reqIndex ? way0V_124 : _GEN_262; // @[DCache.scala 120:{33,33}]
  wire  _GEN_264 = 7'h7d == reqIndex ? way0V_125 : _GEN_263; // @[DCache.scala 120:{33,33}]
  wire  _GEN_265 = 7'h7e == reqIndex ? way0V_126 : _GEN_264; // @[DCache.scala 120:{33,33}]
  wire  _GEN_266 = 7'h7f == reqIndex ? way0V_127 : _GEN_265; // @[DCache.scala 120:{33,33}]
  wire [20:0] _GEN_12 = 7'h1 == reqIndex ? way0Tag_1 : way0Tag_0; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_13 = 7'h2 == reqIndex ? way0Tag_2 : _GEN_12; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_14 = 7'h3 == reqIndex ? way0Tag_3 : _GEN_13; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_15 = 7'h4 == reqIndex ? way0Tag_4 : _GEN_14; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_16 = 7'h5 == reqIndex ? way0Tag_5 : _GEN_15; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_17 = 7'h6 == reqIndex ? way0Tag_6 : _GEN_16; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_18 = 7'h7 == reqIndex ? way0Tag_7 : _GEN_17; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_19 = 7'h8 == reqIndex ? way0Tag_8 : _GEN_18; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_20 = 7'h9 == reqIndex ? way0Tag_9 : _GEN_19; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_21 = 7'ha == reqIndex ? way0Tag_10 : _GEN_20; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_22 = 7'hb == reqIndex ? way0Tag_11 : _GEN_21; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_23 = 7'hc == reqIndex ? way0Tag_12 : _GEN_22; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_24 = 7'hd == reqIndex ? way0Tag_13 : _GEN_23; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_25 = 7'he == reqIndex ? way0Tag_14 : _GEN_24; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_26 = 7'hf == reqIndex ? way0Tag_15 : _GEN_25; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_27 = 7'h10 == reqIndex ? way0Tag_16 : _GEN_26; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_28 = 7'h11 == reqIndex ? way0Tag_17 : _GEN_27; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_29 = 7'h12 == reqIndex ? way0Tag_18 : _GEN_28; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_30 = 7'h13 == reqIndex ? way0Tag_19 : _GEN_29; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_31 = 7'h14 == reqIndex ? way0Tag_20 : _GEN_30; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_32 = 7'h15 == reqIndex ? way0Tag_21 : _GEN_31; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_33 = 7'h16 == reqIndex ? way0Tag_22 : _GEN_32; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_34 = 7'h17 == reqIndex ? way0Tag_23 : _GEN_33; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_35 = 7'h18 == reqIndex ? way0Tag_24 : _GEN_34; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_36 = 7'h19 == reqIndex ? way0Tag_25 : _GEN_35; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_37 = 7'h1a == reqIndex ? way0Tag_26 : _GEN_36; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_38 = 7'h1b == reqIndex ? way0Tag_27 : _GEN_37; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_39 = 7'h1c == reqIndex ? way0Tag_28 : _GEN_38; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_40 = 7'h1d == reqIndex ? way0Tag_29 : _GEN_39; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_41 = 7'h1e == reqIndex ? way0Tag_30 : _GEN_40; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_42 = 7'h1f == reqIndex ? way0Tag_31 : _GEN_41; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_43 = 7'h20 == reqIndex ? way0Tag_32 : _GEN_42; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_44 = 7'h21 == reqIndex ? way0Tag_33 : _GEN_43; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_45 = 7'h22 == reqIndex ? way0Tag_34 : _GEN_44; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_46 = 7'h23 == reqIndex ? way0Tag_35 : _GEN_45; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_47 = 7'h24 == reqIndex ? way0Tag_36 : _GEN_46; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_48 = 7'h25 == reqIndex ? way0Tag_37 : _GEN_47; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_49 = 7'h26 == reqIndex ? way0Tag_38 : _GEN_48; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_50 = 7'h27 == reqIndex ? way0Tag_39 : _GEN_49; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_51 = 7'h28 == reqIndex ? way0Tag_40 : _GEN_50; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_52 = 7'h29 == reqIndex ? way0Tag_41 : _GEN_51; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_53 = 7'h2a == reqIndex ? way0Tag_42 : _GEN_52; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_54 = 7'h2b == reqIndex ? way0Tag_43 : _GEN_53; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_55 = 7'h2c == reqIndex ? way0Tag_44 : _GEN_54; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_56 = 7'h2d == reqIndex ? way0Tag_45 : _GEN_55; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_57 = 7'h2e == reqIndex ? way0Tag_46 : _GEN_56; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_58 = 7'h2f == reqIndex ? way0Tag_47 : _GEN_57; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_59 = 7'h30 == reqIndex ? way0Tag_48 : _GEN_58; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_60 = 7'h31 == reqIndex ? way0Tag_49 : _GEN_59; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_61 = 7'h32 == reqIndex ? way0Tag_50 : _GEN_60; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_62 = 7'h33 == reqIndex ? way0Tag_51 : _GEN_61; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_63 = 7'h34 == reqIndex ? way0Tag_52 : _GEN_62; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_64 = 7'h35 == reqIndex ? way0Tag_53 : _GEN_63; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_65 = 7'h36 == reqIndex ? way0Tag_54 : _GEN_64; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_66 = 7'h37 == reqIndex ? way0Tag_55 : _GEN_65; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_67 = 7'h38 == reqIndex ? way0Tag_56 : _GEN_66; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_68 = 7'h39 == reqIndex ? way0Tag_57 : _GEN_67; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_69 = 7'h3a == reqIndex ? way0Tag_58 : _GEN_68; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_70 = 7'h3b == reqIndex ? way0Tag_59 : _GEN_69; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_71 = 7'h3c == reqIndex ? way0Tag_60 : _GEN_70; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_72 = 7'h3d == reqIndex ? way0Tag_61 : _GEN_71; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_73 = 7'h3e == reqIndex ? way0Tag_62 : _GEN_72; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_74 = 7'h3f == reqIndex ? way0Tag_63 : _GEN_73; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_75 = 7'h40 == reqIndex ? way0Tag_64 : _GEN_74; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_76 = 7'h41 == reqIndex ? way0Tag_65 : _GEN_75; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_77 = 7'h42 == reqIndex ? way0Tag_66 : _GEN_76; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_78 = 7'h43 == reqIndex ? way0Tag_67 : _GEN_77; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_79 = 7'h44 == reqIndex ? way0Tag_68 : _GEN_78; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_80 = 7'h45 == reqIndex ? way0Tag_69 : _GEN_79; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_81 = 7'h46 == reqIndex ? way0Tag_70 : _GEN_80; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_82 = 7'h47 == reqIndex ? way0Tag_71 : _GEN_81; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_83 = 7'h48 == reqIndex ? way0Tag_72 : _GEN_82; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_84 = 7'h49 == reqIndex ? way0Tag_73 : _GEN_83; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_85 = 7'h4a == reqIndex ? way0Tag_74 : _GEN_84; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_86 = 7'h4b == reqIndex ? way0Tag_75 : _GEN_85; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_87 = 7'h4c == reqIndex ? way0Tag_76 : _GEN_86; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_88 = 7'h4d == reqIndex ? way0Tag_77 : _GEN_87; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_89 = 7'h4e == reqIndex ? way0Tag_78 : _GEN_88; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_90 = 7'h4f == reqIndex ? way0Tag_79 : _GEN_89; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_91 = 7'h50 == reqIndex ? way0Tag_80 : _GEN_90; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_92 = 7'h51 == reqIndex ? way0Tag_81 : _GEN_91; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_93 = 7'h52 == reqIndex ? way0Tag_82 : _GEN_92; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_94 = 7'h53 == reqIndex ? way0Tag_83 : _GEN_93; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_95 = 7'h54 == reqIndex ? way0Tag_84 : _GEN_94; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_96 = 7'h55 == reqIndex ? way0Tag_85 : _GEN_95; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_97 = 7'h56 == reqIndex ? way0Tag_86 : _GEN_96; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_98 = 7'h57 == reqIndex ? way0Tag_87 : _GEN_97; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_99 = 7'h58 == reqIndex ? way0Tag_88 : _GEN_98; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_100 = 7'h59 == reqIndex ? way0Tag_89 : _GEN_99; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_101 = 7'h5a == reqIndex ? way0Tag_90 : _GEN_100; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_102 = 7'h5b == reqIndex ? way0Tag_91 : _GEN_101; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_103 = 7'h5c == reqIndex ? way0Tag_92 : _GEN_102; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_104 = 7'h5d == reqIndex ? way0Tag_93 : _GEN_103; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_105 = 7'h5e == reqIndex ? way0Tag_94 : _GEN_104; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_106 = 7'h5f == reqIndex ? way0Tag_95 : _GEN_105; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_107 = 7'h60 == reqIndex ? way0Tag_96 : _GEN_106; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_108 = 7'h61 == reqIndex ? way0Tag_97 : _GEN_107; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_109 = 7'h62 == reqIndex ? way0Tag_98 : _GEN_108; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_110 = 7'h63 == reqIndex ? way0Tag_99 : _GEN_109; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_111 = 7'h64 == reqIndex ? way0Tag_100 : _GEN_110; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_112 = 7'h65 == reqIndex ? way0Tag_101 : _GEN_111; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_113 = 7'h66 == reqIndex ? way0Tag_102 : _GEN_112; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_114 = 7'h67 == reqIndex ? way0Tag_103 : _GEN_113; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_115 = 7'h68 == reqIndex ? way0Tag_104 : _GEN_114; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_116 = 7'h69 == reqIndex ? way0Tag_105 : _GEN_115; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_117 = 7'h6a == reqIndex ? way0Tag_106 : _GEN_116; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_118 = 7'h6b == reqIndex ? way0Tag_107 : _GEN_117; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_119 = 7'h6c == reqIndex ? way0Tag_108 : _GEN_118; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_120 = 7'h6d == reqIndex ? way0Tag_109 : _GEN_119; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_121 = 7'h6e == reqIndex ? way0Tag_110 : _GEN_120; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_122 = 7'h6f == reqIndex ? way0Tag_111 : _GEN_121; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_123 = 7'h70 == reqIndex ? way0Tag_112 : _GEN_122; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_124 = 7'h71 == reqIndex ? way0Tag_113 : _GEN_123; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_125 = 7'h72 == reqIndex ? way0Tag_114 : _GEN_124; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_126 = 7'h73 == reqIndex ? way0Tag_115 : _GEN_125; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_127 = 7'h74 == reqIndex ? way0Tag_116 : _GEN_126; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_128 = 7'h75 == reqIndex ? way0Tag_117 : _GEN_127; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_129 = 7'h76 == reqIndex ? way0Tag_118 : _GEN_128; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_130 = 7'h77 == reqIndex ? way0Tag_119 : _GEN_129; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_131 = 7'h78 == reqIndex ? way0Tag_120 : _GEN_130; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_132 = 7'h79 == reqIndex ? way0Tag_121 : _GEN_131; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_133 = 7'h7a == reqIndex ? way0Tag_122 : _GEN_132; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_134 = 7'h7b == reqIndex ? way0Tag_123 : _GEN_133; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_135 = 7'h7c == reqIndex ? way0Tag_124 : _GEN_134; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_136 = 7'h7d == reqIndex ? way0Tag_125 : _GEN_135; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_137 = 7'h7e == reqIndex ? way0Tag_126 : _GEN_136; // @[DCache.scala 120:{55,55}]
  wire [20:0] _GEN_138 = 7'h7f == reqIndex ? way0Tag_127 : _GEN_137; // @[DCache.scala 120:{55,55}]
  wire  sHitEn = state == 3'h1; // @[DCache.scala 119:22]
  wire  way0Hit = _GEN_266 & _GEN_138 == reqTag & sHitEn; // @[DCache.scala 120:67]
  wire  _GEN_396 = 7'h1 == reqIndex ? way1V_1 : way1V_0; // @[DCache.scala 121:{33,33}]
  wire  _GEN_397 = 7'h2 == reqIndex ? way1V_2 : _GEN_396; // @[DCache.scala 121:{33,33}]
  wire  _GEN_398 = 7'h3 == reqIndex ? way1V_3 : _GEN_397; // @[DCache.scala 121:{33,33}]
  wire  _GEN_399 = 7'h4 == reqIndex ? way1V_4 : _GEN_398; // @[DCache.scala 121:{33,33}]
  wire  _GEN_400 = 7'h5 == reqIndex ? way1V_5 : _GEN_399; // @[DCache.scala 121:{33,33}]
  wire  _GEN_401 = 7'h6 == reqIndex ? way1V_6 : _GEN_400; // @[DCache.scala 121:{33,33}]
  wire  _GEN_402 = 7'h7 == reqIndex ? way1V_7 : _GEN_401; // @[DCache.scala 121:{33,33}]
  wire  _GEN_403 = 7'h8 == reqIndex ? way1V_8 : _GEN_402; // @[DCache.scala 121:{33,33}]
  wire  _GEN_404 = 7'h9 == reqIndex ? way1V_9 : _GEN_403; // @[DCache.scala 121:{33,33}]
  wire  _GEN_405 = 7'ha == reqIndex ? way1V_10 : _GEN_404; // @[DCache.scala 121:{33,33}]
  wire  _GEN_406 = 7'hb == reqIndex ? way1V_11 : _GEN_405; // @[DCache.scala 121:{33,33}]
  wire  _GEN_407 = 7'hc == reqIndex ? way1V_12 : _GEN_406; // @[DCache.scala 121:{33,33}]
  wire  _GEN_408 = 7'hd == reqIndex ? way1V_13 : _GEN_407; // @[DCache.scala 121:{33,33}]
  wire  _GEN_409 = 7'he == reqIndex ? way1V_14 : _GEN_408; // @[DCache.scala 121:{33,33}]
  wire  _GEN_410 = 7'hf == reqIndex ? way1V_15 : _GEN_409; // @[DCache.scala 121:{33,33}]
  wire  _GEN_411 = 7'h10 == reqIndex ? way1V_16 : _GEN_410; // @[DCache.scala 121:{33,33}]
  wire  _GEN_412 = 7'h11 == reqIndex ? way1V_17 : _GEN_411; // @[DCache.scala 121:{33,33}]
  wire  _GEN_413 = 7'h12 == reqIndex ? way1V_18 : _GEN_412; // @[DCache.scala 121:{33,33}]
  wire  _GEN_414 = 7'h13 == reqIndex ? way1V_19 : _GEN_413; // @[DCache.scala 121:{33,33}]
  wire  _GEN_415 = 7'h14 == reqIndex ? way1V_20 : _GEN_414; // @[DCache.scala 121:{33,33}]
  wire  _GEN_416 = 7'h15 == reqIndex ? way1V_21 : _GEN_415; // @[DCache.scala 121:{33,33}]
  wire  _GEN_417 = 7'h16 == reqIndex ? way1V_22 : _GEN_416; // @[DCache.scala 121:{33,33}]
  wire  _GEN_418 = 7'h17 == reqIndex ? way1V_23 : _GEN_417; // @[DCache.scala 121:{33,33}]
  wire  _GEN_419 = 7'h18 == reqIndex ? way1V_24 : _GEN_418; // @[DCache.scala 121:{33,33}]
  wire  _GEN_420 = 7'h19 == reqIndex ? way1V_25 : _GEN_419; // @[DCache.scala 121:{33,33}]
  wire  _GEN_421 = 7'h1a == reqIndex ? way1V_26 : _GEN_420; // @[DCache.scala 121:{33,33}]
  wire  _GEN_422 = 7'h1b == reqIndex ? way1V_27 : _GEN_421; // @[DCache.scala 121:{33,33}]
  wire  _GEN_423 = 7'h1c == reqIndex ? way1V_28 : _GEN_422; // @[DCache.scala 121:{33,33}]
  wire  _GEN_424 = 7'h1d == reqIndex ? way1V_29 : _GEN_423; // @[DCache.scala 121:{33,33}]
  wire  _GEN_425 = 7'h1e == reqIndex ? way1V_30 : _GEN_424; // @[DCache.scala 121:{33,33}]
  wire  _GEN_426 = 7'h1f == reqIndex ? way1V_31 : _GEN_425; // @[DCache.scala 121:{33,33}]
  wire  _GEN_427 = 7'h20 == reqIndex ? way1V_32 : _GEN_426; // @[DCache.scala 121:{33,33}]
  wire  _GEN_428 = 7'h21 == reqIndex ? way1V_33 : _GEN_427; // @[DCache.scala 121:{33,33}]
  wire  _GEN_429 = 7'h22 == reqIndex ? way1V_34 : _GEN_428; // @[DCache.scala 121:{33,33}]
  wire  _GEN_430 = 7'h23 == reqIndex ? way1V_35 : _GEN_429; // @[DCache.scala 121:{33,33}]
  wire  _GEN_431 = 7'h24 == reqIndex ? way1V_36 : _GEN_430; // @[DCache.scala 121:{33,33}]
  wire  _GEN_432 = 7'h25 == reqIndex ? way1V_37 : _GEN_431; // @[DCache.scala 121:{33,33}]
  wire  _GEN_433 = 7'h26 == reqIndex ? way1V_38 : _GEN_432; // @[DCache.scala 121:{33,33}]
  wire  _GEN_434 = 7'h27 == reqIndex ? way1V_39 : _GEN_433; // @[DCache.scala 121:{33,33}]
  wire  _GEN_435 = 7'h28 == reqIndex ? way1V_40 : _GEN_434; // @[DCache.scala 121:{33,33}]
  wire  _GEN_436 = 7'h29 == reqIndex ? way1V_41 : _GEN_435; // @[DCache.scala 121:{33,33}]
  wire  _GEN_437 = 7'h2a == reqIndex ? way1V_42 : _GEN_436; // @[DCache.scala 121:{33,33}]
  wire  _GEN_438 = 7'h2b == reqIndex ? way1V_43 : _GEN_437; // @[DCache.scala 121:{33,33}]
  wire  _GEN_439 = 7'h2c == reqIndex ? way1V_44 : _GEN_438; // @[DCache.scala 121:{33,33}]
  wire  _GEN_440 = 7'h2d == reqIndex ? way1V_45 : _GEN_439; // @[DCache.scala 121:{33,33}]
  wire  _GEN_441 = 7'h2e == reqIndex ? way1V_46 : _GEN_440; // @[DCache.scala 121:{33,33}]
  wire  _GEN_442 = 7'h2f == reqIndex ? way1V_47 : _GEN_441; // @[DCache.scala 121:{33,33}]
  wire  _GEN_443 = 7'h30 == reqIndex ? way1V_48 : _GEN_442; // @[DCache.scala 121:{33,33}]
  wire  _GEN_444 = 7'h31 == reqIndex ? way1V_49 : _GEN_443; // @[DCache.scala 121:{33,33}]
  wire  _GEN_445 = 7'h32 == reqIndex ? way1V_50 : _GEN_444; // @[DCache.scala 121:{33,33}]
  wire  _GEN_446 = 7'h33 == reqIndex ? way1V_51 : _GEN_445; // @[DCache.scala 121:{33,33}]
  wire  _GEN_447 = 7'h34 == reqIndex ? way1V_52 : _GEN_446; // @[DCache.scala 121:{33,33}]
  wire  _GEN_448 = 7'h35 == reqIndex ? way1V_53 : _GEN_447; // @[DCache.scala 121:{33,33}]
  wire  _GEN_449 = 7'h36 == reqIndex ? way1V_54 : _GEN_448; // @[DCache.scala 121:{33,33}]
  wire  _GEN_450 = 7'h37 == reqIndex ? way1V_55 : _GEN_449; // @[DCache.scala 121:{33,33}]
  wire  _GEN_451 = 7'h38 == reqIndex ? way1V_56 : _GEN_450; // @[DCache.scala 121:{33,33}]
  wire  _GEN_452 = 7'h39 == reqIndex ? way1V_57 : _GEN_451; // @[DCache.scala 121:{33,33}]
  wire  _GEN_453 = 7'h3a == reqIndex ? way1V_58 : _GEN_452; // @[DCache.scala 121:{33,33}]
  wire  _GEN_454 = 7'h3b == reqIndex ? way1V_59 : _GEN_453; // @[DCache.scala 121:{33,33}]
  wire  _GEN_455 = 7'h3c == reqIndex ? way1V_60 : _GEN_454; // @[DCache.scala 121:{33,33}]
  wire  _GEN_456 = 7'h3d == reqIndex ? way1V_61 : _GEN_455; // @[DCache.scala 121:{33,33}]
  wire  _GEN_457 = 7'h3e == reqIndex ? way1V_62 : _GEN_456; // @[DCache.scala 121:{33,33}]
  wire  _GEN_458 = 7'h3f == reqIndex ? way1V_63 : _GEN_457; // @[DCache.scala 121:{33,33}]
  wire  _GEN_459 = 7'h40 == reqIndex ? way1V_64 : _GEN_458; // @[DCache.scala 121:{33,33}]
  wire  _GEN_460 = 7'h41 == reqIndex ? way1V_65 : _GEN_459; // @[DCache.scala 121:{33,33}]
  wire  _GEN_461 = 7'h42 == reqIndex ? way1V_66 : _GEN_460; // @[DCache.scala 121:{33,33}]
  wire  _GEN_462 = 7'h43 == reqIndex ? way1V_67 : _GEN_461; // @[DCache.scala 121:{33,33}]
  wire  _GEN_463 = 7'h44 == reqIndex ? way1V_68 : _GEN_462; // @[DCache.scala 121:{33,33}]
  wire  _GEN_464 = 7'h45 == reqIndex ? way1V_69 : _GEN_463; // @[DCache.scala 121:{33,33}]
  wire  _GEN_465 = 7'h46 == reqIndex ? way1V_70 : _GEN_464; // @[DCache.scala 121:{33,33}]
  wire  _GEN_466 = 7'h47 == reqIndex ? way1V_71 : _GEN_465; // @[DCache.scala 121:{33,33}]
  wire  _GEN_467 = 7'h48 == reqIndex ? way1V_72 : _GEN_466; // @[DCache.scala 121:{33,33}]
  wire  _GEN_468 = 7'h49 == reqIndex ? way1V_73 : _GEN_467; // @[DCache.scala 121:{33,33}]
  wire  _GEN_469 = 7'h4a == reqIndex ? way1V_74 : _GEN_468; // @[DCache.scala 121:{33,33}]
  wire  _GEN_470 = 7'h4b == reqIndex ? way1V_75 : _GEN_469; // @[DCache.scala 121:{33,33}]
  wire  _GEN_471 = 7'h4c == reqIndex ? way1V_76 : _GEN_470; // @[DCache.scala 121:{33,33}]
  wire  _GEN_472 = 7'h4d == reqIndex ? way1V_77 : _GEN_471; // @[DCache.scala 121:{33,33}]
  wire  _GEN_473 = 7'h4e == reqIndex ? way1V_78 : _GEN_472; // @[DCache.scala 121:{33,33}]
  wire  _GEN_474 = 7'h4f == reqIndex ? way1V_79 : _GEN_473; // @[DCache.scala 121:{33,33}]
  wire  _GEN_475 = 7'h50 == reqIndex ? way1V_80 : _GEN_474; // @[DCache.scala 121:{33,33}]
  wire  _GEN_476 = 7'h51 == reqIndex ? way1V_81 : _GEN_475; // @[DCache.scala 121:{33,33}]
  wire  _GEN_477 = 7'h52 == reqIndex ? way1V_82 : _GEN_476; // @[DCache.scala 121:{33,33}]
  wire  _GEN_478 = 7'h53 == reqIndex ? way1V_83 : _GEN_477; // @[DCache.scala 121:{33,33}]
  wire  _GEN_479 = 7'h54 == reqIndex ? way1V_84 : _GEN_478; // @[DCache.scala 121:{33,33}]
  wire  _GEN_480 = 7'h55 == reqIndex ? way1V_85 : _GEN_479; // @[DCache.scala 121:{33,33}]
  wire  _GEN_481 = 7'h56 == reqIndex ? way1V_86 : _GEN_480; // @[DCache.scala 121:{33,33}]
  wire  _GEN_482 = 7'h57 == reqIndex ? way1V_87 : _GEN_481; // @[DCache.scala 121:{33,33}]
  wire  _GEN_483 = 7'h58 == reqIndex ? way1V_88 : _GEN_482; // @[DCache.scala 121:{33,33}]
  wire  _GEN_484 = 7'h59 == reqIndex ? way1V_89 : _GEN_483; // @[DCache.scala 121:{33,33}]
  wire  _GEN_485 = 7'h5a == reqIndex ? way1V_90 : _GEN_484; // @[DCache.scala 121:{33,33}]
  wire  _GEN_486 = 7'h5b == reqIndex ? way1V_91 : _GEN_485; // @[DCache.scala 121:{33,33}]
  wire  _GEN_487 = 7'h5c == reqIndex ? way1V_92 : _GEN_486; // @[DCache.scala 121:{33,33}]
  wire  _GEN_488 = 7'h5d == reqIndex ? way1V_93 : _GEN_487; // @[DCache.scala 121:{33,33}]
  wire  _GEN_489 = 7'h5e == reqIndex ? way1V_94 : _GEN_488; // @[DCache.scala 121:{33,33}]
  wire  _GEN_490 = 7'h5f == reqIndex ? way1V_95 : _GEN_489; // @[DCache.scala 121:{33,33}]
  wire  _GEN_491 = 7'h60 == reqIndex ? way1V_96 : _GEN_490; // @[DCache.scala 121:{33,33}]
  wire  _GEN_492 = 7'h61 == reqIndex ? way1V_97 : _GEN_491; // @[DCache.scala 121:{33,33}]
  wire  _GEN_493 = 7'h62 == reqIndex ? way1V_98 : _GEN_492; // @[DCache.scala 121:{33,33}]
  wire  _GEN_494 = 7'h63 == reqIndex ? way1V_99 : _GEN_493; // @[DCache.scala 121:{33,33}]
  wire  _GEN_495 = 7'h64 == reqIndex ? way1V_100 : _GEN_494; // @[DCache.scala 121:{33,33}]
  wire  _GEN_496 = 7'h65 == reqIndex ? way1V_101 : _GEN_495; // @[DCache.scala 121:{33,33}]
  wire  _GEN_497 = 7'h66 == reqIndex ? way1V_102 : _GEN_496; // @[DCache.scala 121:{33,33}]
  wire  _GEN_498 = 7'h67 == reqIndex ? way1V_103 : _GEN_497; // @[DCache.scala 121:{33,33}]
  wire  _GEN_499 = 7'h68 == reqIndex ? way1V_104 : _GEN_498; // @[DCache.scala 121:{33,33}]
  wire  _GEN_500 = 7'h69 == reqIndex ? way1V_105 : _GEN_499; // @[DCache.scala 121:{33,33}]
  wire  _GEN_501 = 7'h6a == reqIndex ? way1V_106 : _GEN_500; // @[DCache.scala 121:{33,33}]
  wire  _GEN_502 = 7'h6b == reqIndex ? way1V_107 : _GEN_501; // @[DCache.scala 121:{33,33}]
  wire  _GEN_503 = 7'h6c == reqIndex ? way1V_108 : _GEN_502; // @[DCache.scala 121:{33,33}]
  wire  _GEN_504 = 7'h6d == reqIndex ? way1V_109 : _GEN_503; // @[DCache.scala 121:{33,33}]
  wire  _GEN_505 = 7'h6e == reqIndex ? way1V_110 : _GEN_504; // @[DCache.scala 121:{33,33}]
  wire  _GEN_506 = 7'h6f == reqIndex ? way1V_111 : _GEN_505; // @[DCache.scala 121:{33,33}]
  wire  _GEN_507 = 7'h70 == reqIndex ? way1V_112 : _GEN_506; // @[DCache.scala 121:{33,33}]
  wire  _GEN_508 = 7'h71 == reqIndex ? way1V_113 : _GEN_507; // @[DCache.scala 121:{33,33}]
  wire  _GEN_509 = 7'h72 == reqIndex ? way1V_114 : _GEN_508; // @[DCache.scala 121:{33,33}]
  wire  _GEN_510 = 7'h73 == reqIndex ? way1V_115 : _GEN_509; // @[DCache.scala 121:{33,33}]
  wire  _GEN_511 = 7'h74 == reqIndex ? way1V_116 : _GEN_510; // @[DCache.scala 121:{33,33}]
  wire  _GEN_512 = 7'h75 == reqIndex ? way1V_117 : _GEN_511; // @[DCache.scala 121:{33,33}]
  wire  _GEN_513 = 7'h76 == reqIndex ? way1V_118 : _GEN_512; // @[DCache.scala 121:{33,33}]
  wire  _GEN_514 = 7'h77 == reqIndex ? way1V_119 : _GEN_513; // @[DCache.scala 121:{33,33}]
  wire  _GEN_515 = 7'h78 == reqIndex ? way1V_120 : _GEN_514; // @[DCache.scala 121:{33,33}]
  wire  _GEN_516 = 7'h79 == reqIndex ? way1V_121 : _GEN_515; // @[DCache.scala 121:{33,33}]
  wire  _GEN_517 = 7'h7a == reqIndex ? way1V_122 : _GEN_516; // @[DCache.scala 121:{33,33}]
  wire  _GEN_518 = 7'h7b == reqIndex ? way1V_123 : _GEN_517; // @[DCache.scala 121:{33,33}]
  wire  _GEN_519 = 7'h7c == reqIndex ? way1V_124 : _GEN_518; // @[DCache.scala 121:{33,33}]
  wire  _GEN_520 = 7'h7d == reqIndex ? way1V_125 : _GEN_519; // @[DCache.scala 121:{33,33}]
  wire  _GEN_521 = 7'h7e == reqIndex ? way1V_126 : _GEN_520; // @[DCache.scala 121:{33,33}]
  wire  _GEN_522 = 7'h7f == reqIndex ? way1V_127 : _GEN_521; // @[DCache.scala 121:{33,33}]
  wire [20:0] _GEN_268 = 7'h1 == reqIndex ? way1Tag_1 : way1Tag_0; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_269 = 7'h2 == reqIndex ? way1Tag_2 : _GEN_268; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_270 = 7'h3 == reqIndex ? way1Tag_3 : _GEN_269; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_271 = 7'h4 == reqIndex ? way1Tag_4 : _GEN_270; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_272 = 7'h5 == reqIndex ? way1Tag_5 : _GEN_271; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_273 = 7'h6 == reqIndex ? way1Tag_6 : _GEN_272; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_274 = 7'h7 == reqIndex ? way1Tag_7 : _GEN_273; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_275 = 7'h8 == reqIndex ? way1Tag_8 : _GEN_274; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_276 = 7'h9 == reqIndex ? way1Tag_9 : _GEN_275; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_277 = 7'ha == reqIndex ? way1Tag_10 : _GEN_276; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_278 = 7'hb == reqIndex ? way1Tag_11 : _GEN_277; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_279 = 7'hc == reqIndex ? way1Tag_12 : _GEN_278; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_280 = 7'hd == reqIndex ? way1Tag_13 : _GEN_279; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_281 = 7'he == reqIndex ? way1Tag_14 : _GEN_280; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_282 = 7'hf == reqIndex ? way1Tag_15 : _GEN_281; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_283 = 7'h10 == reqIndex ? way1Tag_16 : _GEN_282; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_284 = 7'h11 == reqIndex ? way1Tag_17 : _GEN_283; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_285 = 7'h12 == reqIndex ? way1Tag_18 : _GEN_284; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_286 = 7'h13 == reqIndex ? way1Tag_19 : _GEN_285; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_287 = 7'h14 == reqIndex ? way1Tag_20 : _GEN_286; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_288 = 7'h15 == reqIndex ? way1Tag_21 : _GEN_287; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_289 = 7'h16 == reqIndex ? way1Tag_22 : _GEN_288; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_290 = 7'h17 == reqIndex ? way1Tag_23 : _GEN_289; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_291 = 7'h18 == reqIndex ? way1Tag_24 : _GEN_290; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_292 = 7'h19 == reqIndex ? way1Tag_25 : _GEN_291; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_293 = 7'h1a == reqIndex ? way1Tag_26 : _GEN_292; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_294 = 7'h1b == reqIndex ? way1Tag_27 : _GEN_293; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_295 = 7'h1c == reqIndex ? way1Tag_28 : _GEN_294; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_296 = 7'h1d == reqIndex ? way1Tag_29 : _GEN_295; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_297 = 7'h1e == reqIndex ? way1Tag_30 : _GEN_296; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_298 = 7'h1f == reqIndex ? way1Tag_31 : _GEN_297; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_299 = 7'h20 == reqIndex ? way1Tag_32 : _GEN_298; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_300 = 7'h21 == reqIndex ? way1Tag_33 : _GEN_299; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_301 = 7'h22 == reqIndex ? way1Tag_34 : _GEN_300; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_302 = 7'h23 == reqIndex ? way1Tag_35 : _GEN_301; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_303 = 7'h24 == reqIndex ? way1Tag_36 : _GEN_302; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_304 = 7'h25 == reqIndex ? way1Tag_37 : _GEN_303; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_305 = 7'h26 == reqIndex ? way1Tag_38 : _GEN_304; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_306 = 7'h27 == reqIndex ? way1Tag_39 : _GEN_305; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_307 = 7'h28 == reqIndex ? way1Tag_40 : _GEN_306; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_308 = 7'h29 == reqIndex ? way1Tag_41 : _GEN_307; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_309 = 7'h2a == reqIndex ? way1Tag_42 : _GEN_308; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_310 = 7'h2b == reqIndex ? way1Tag_43 : _GEN_309; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_311 = 7'h2c == reqIndex ? way1Tag_44 : _GEN_310; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_312 = 7'h2d == reqIndex ? way1Tag_45 : _GEN_311; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_313 = 7'h2e == reqIndex ? way1Tag_46 : _GEN_312; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_314 = 7'h2f == reqIndex ? way1Tag_47 : _GEN_313; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_315 = 7'h30 == reqIndex ? way1Tag_48 : _GEN_314; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_316 = 7'h31 == reqIndex ? way1Tag_49 : _GEN_315; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_317 = 7'h32 == reqIndex ? way1Tag_50 : _GEN_316; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_318 = 7'h33 == reqIndex ? way1Tag_51 : _GEN_317; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_319 = 7'h34 == reqIndex ? way1Tag_52 : _GEN_318; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_320 = 7'h35 == reqIndex ? way1Tag_53 : _GEN_319; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_321 = 7'h36 == reqIndex ? way1Tag_54 : _GEN_320; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_322 = 7'h37 == reqIndex ? way1Tag_55 : _GEN_321; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_323 = 7'h38 == reqIndex ? way1Tag_56 : _GEN_322; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_324 = 7'h39 == reqIndex ? way1Tag_57 : _GEN_323; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_325 = 7'h3a == reqIndex ? way1Tag_58 : _GEN_324; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_326 = 7'h3b == reqIndex ? way1Tag_59 : _GEN_325; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_327 = 7'h3c == reqIndex ? way1Tag_60 : _GEN_326; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_328 = 7'h3d == reqIndex ? way1Tag_61 : _GEN_327; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_329 = 7'h3e == reqIndex ? way1Tag_62 : _GEN_328; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_330 = 7'h3f == reqIndex ? way1Tag_63 : _GEN_329; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_331 = 7'h40 == reqIndex ? way1Tag_64 : _GEN_330; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_332 = 7'h41 == reqIndex ? way1Tag_65 : _GEN_331; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_333 = 7'h42 == reqIndex ? way1Tag_66 : _GEN_332; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_334 = 7'h43 == reqIndex ? way1Tag_67 : _GEN_333; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_335 = 7'h44 == reqIndex ? way1Tag_68 : _GEN_334; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_336 = 7'h45 == reqIndex ? way1Tag_69 : _GEN_335; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_337 = 7'h46 == reqIndex ? way1Tag_70 : _GEN_336; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_338 = 7'h47 == reqIndex ? way1Tag_71 : _GEN_337; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_339 = 7'h48 == reqIndex ? way1Tag_72 : _GEN_338; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_340 = 7'h49 == reqIndex ? way1Tag_73 : _GEN_339; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_341 = 7'h4a == reqIndex ? way1Tag_74 : _GEN_340; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_342 = 7'h4b == reqIndex ? way1Tag_75 : _GEN_341; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_343 = 7'h4c == reqIndex ? way1Tag_76 : _GEN_342; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_344 = 7'h4d == reqIndex ? way1Tag_77 : _GEN_343; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_345 = 7'h4e == reqIndex ? way1Tag_78 : _GEN_344; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_346 = 7'h4f == reqIndex ? way1Tag_79 : _GEN_345; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_347 = 7'h50 == reqIndex ? way1Tag_80 : _GEN_346; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_348 = 7'h51 == reqIndex ? way1Tag_81 : _GEN_347; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_349 = 7'h52 == reqIndex ? way1Tag_82 : _GEN_348; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_350 = 7'h53 == reqIndex ? way1Tag_83 : _GEN_349; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_351 = 7'h54 == reqIndex ? way1Tag_84 : _GEN_350; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_352 = 7'h55 == reqIndex ? way1Tag_85 : _GEN_351; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_353 = 7'h56 == reqIndex ? way1Tag_86 : _GEN_352; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_354 = 7'h57 == reqIndex ? way1Tag_87 : _GEN_353; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_355 = 7'h58 == reqIndex ? way1Tag_88 : _GEN_354; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_356 = 7'h59 == reqIndex ? way1Tag_89 : _GEN_355; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_357 = 7'h5a == reqIndex ? way1Tag_90 : _GEN_356; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_358 = 7'h5b == reqIndex ? way1Tag_91 : _GEN_357; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_359 = 7'h5c == reqIndex ? way1Tag_92 : _GEN_358; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_360 = 7'h5d == reqIndex ? way1Tag_93 : _GEN_359; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_361 = 7'h5e == reqIndex ? way1Tag_94 : _GEN_360; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_362 = 7'h5f == reqIndex ? way1Tag_95 : _GEN_361; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_363 = 7'h60 == reqIndex ? way1Tag_96 : _GEN_362; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_364 = 7'h61 == reqIndex ? way1Tag_97 : _GEN_363; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_365 = 7'h62 == reqIndex ? way1Tag_98 : _GEN_364; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_366 = 7'h63 == reqIndex ? way1Tag_99 : _GEN_365; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_367 = 7'h64 == reqIndex ? way1Tag_100 : _GEN_366; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_368 = 7'h65 == reqIndex ? way1Tag_101 : _GEN_367; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_369 = 7'h66 == reqIndex ? way1Tag_102 : _GEN_368; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_370 = 7'h67 == reqIndex ? way1Tag_103 : _GEN_369; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_371 = 7'h68 == reqIndex ? way1Tag_104 : _GEN_370; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_372 = 7'h69 == reqIndex ? way1Tag_105 : _GEN_371; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_373 = 7'h6a == reqIndex ? way1Tag_106 : _GEN_372; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_374 = 7'h6b == reqIndex ? way1Tag_107 : _GEN_373; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_375 = 7'h6c == reqIndex ? way1Tag_108 : _GEN_374; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_376 = 7'h6d == reqIndex ? way1Tag_109 : _GEN_375; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_377 = 7'h6e == reqIndex ? way1Tag_110 : _GEN_376; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_378 = 7'h6f == reqIndex ? way1Tag_111 : _GEN_377; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_379 = 7'h70 == reqIndex ? way1Tag_112 : _GEN_378; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_380 = 7'h71 == reqIndex ? way1Tag_113 : _GEN_379; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_381 = 7'h72 == reqIndex ? way1Tag_114 : _GEN_380; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_382 = 7'h73 == reqIndex ? way1Tag_115 : _GEN_381; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_383 = 7'h74 == reqIndex ? way1Tag_116 : _GEN_382; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_384 = 7'h75 == reqIndex ? way1Tag_117 : _GEN_383; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_385 = 7'h76 == reqIndex ? way1Tag_118 : _GEN_384; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_386 = 7'h77 == reqIndex ? way1Tag_119 : _GEN_385; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_387 = 7'h78 == reqIndex ? way1Tag_120 : _GEN_386; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_388 = 7'h79 == reqIndex ? way1Tag_121 : _GEN_387; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_389 = 7'h7a == reqIndex ? way1Tag_122 : _GEN_388; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_390 = 7'h7b == reqIndex ? way1Tag_123 : _GEN_389; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_391 = 7'h7c == reqIndex ? way1Tag_124 : _GEN_390; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_392 = 7'h7d == reqIndex ? way1Tag_125 : _GEN_391; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_393 = 7'h7e == reqIndex ? way1Tag_126 : _GEN_392; // @[DCache.scala 121:{55,55}]
  wire [20:0] _GEN_394 = 7'h7f == reqIndex ? way1Tag_127 : _GEN_393; // @[DCache.scala 121:{55,55}]
  wire  way1Hit = _GEN_522 & _GEN_394 == reqTag & sHitEn; // @[DCache.scala 121:67]
  wire  cacheHitEn = (way0Hit | way1Hit) & sHitEn; // @[DCache.scala 122:39]
  wire  _GEN_524 = 7'h1 == reqIndex ? way0Age_1 : way0Age_0; // @[DCache.scala 125:{53,53}]
  wire  _GEN_525 = 7'h2 == reqIndex ? way0Age_2 : _GEN_524; // @[DCache.scala 125:{53,53}]
  wire  _GEN_526 = 7'h3 == reqIndex ? way0Age_3 : _GEN_525; // @[DCache.scala 125:{53,53}]
  wire  _GEN_527 = 7'h4 == reqIndex ? way0Age_4 : _GEN_526; // @[DCache.scala 125:{53,53}]
  wire  _GEN_528 = 7'h5 == reqIndex ? way0Age_5 : _GEN_527; // @[DCache.scala 125:{53,53}]
  wire  _GEN_529 = 7'h6 == reqIndex ? way0Age_6 : _GEN_528; // @[DCache.scala 125:{53,53}]
  wire  _GEN_530 = 7'h7 == reqIndex ? way0Age_7 : _GEN_529; // @[DCache.scala 125:{53,53}]
  wire  _GEN_531 = 7'h8 == reqIndex ? way0Age_8 : _GEN_530; // @[DCache.scala 125:{53,53}]
  wire  _GEN_532 = 7'h9 == reqIndex ? way0Age_9 : _GEN_531; // @[DCache.scala 125:{53,53}]
  wire  _GEN_533 = 7'ha == reqIndex ? way0Age_10 : _GEN_532; // @[DCache.scala 125:{53,53}]
  wire  _GEN_534 = 7'hb == reqIndex ? way0Age_11 : _GEN_533; // @[DCache.scala 125:{53,53}]
  wire  _GEN_535 = 7'hc == reqIndex ? way0Age_12 : _GEN_534; // @[DCache.scala 125:{53,53}]
  wire  _GEN_536 = 7'hd == reqIndex ? way0Age_13 : _GEN_535; // @[DCache.scala 125:{53,53}]
  wire  _GEN_537 = 7'he == reqIndex ? way0Age_14 : _GEN_536; // @[DCache.scala 125:{53,53}]
  wire  _GEN_538 = 7'hf == reqIndex ? way0Age_15 : _GEN_537; // @[DCache.scala 125:{53,53}]
  wire  _GEN_539 = 7'h10 == reqIndex ? way0Age_16 : _GEN_538; // @[DCache.scala 125:{53,53}]
  wire  _GEN_540 = 7'h11 == reqIndex ? way0Age_17 : _GEN_539; // @[DCache.scala 125:{53,53}]
  wire  _GEN_541 = 7'h12 == reqIndex ? way0Age_18 : _GEN_540; // @[DCache.scala 125:{53,53}]
  wire  _GEN_542 = 7'h13 == reqIndex ? way0Age_19 : _GEN_541; // @[DCache.scala 125:{53,53}]
  wire  _GEN_543 = 7'h14 == reqIndex ? way0Age_20 : _GEN_542; // @[DCache.scala 125:{53,53}]
  wire  _GEN_544 = 7'h15 == reqIndex ? way0Age_21 : _GEN_543; // @[DCache.scala 125:{53,53}]
  wire  _GEN_545 = 7'h16 == reqIndex ? way0Age_22 : _GEN_544; // @[DCache.scala 125:{53,53}]
  wire  _GEN_546 = 7'h17 == reqIndex ? way0Age_23 : _GEN_545; // @[DCache.scala 125:{53,53}]
  wire  _GEN_547 = 7'h18 == reqIndex ? way0Age_24 : _GEN_546; // @[DCache.scala 125:{53,53}]
  wire  _GEN_548 = 7'h19 == reqIndex ? way0Age_25 : _GEN_547; // @[DCache.scala 125:{53,53}]
  wire  _GEN_549 = 7'h1a == reqIndex ? way0Age_26 : _GEN_548; // @[DCache.scala 125:{53,53}]
  wire  _GEN_550 = 7'h1b == reqIndex ? way0Age_27 : _GEN_549; // @[DCache.scala 125:{53,53}]
  wire  _GEN_551 = 7'h1c == reqIndex ? way0Age_28 : _GEN_550; // @[DCache.scala 125:{53,53}]
  wire  _GEN_552 = 7'h1d == reqIndex ? way0Age_29 : _GEN_551; // @[DCache.scala 125:{53,53}]
  wire  _GEN_553 = 7'h1e == reqIndex ? way0Age_30 : _GEN_552; // @[DCache.scala 125:{53,53}]
  wire  _GEN_554 = 7'h1f == reqIndex ? way0Age_31 : _GEN_553; // @[DCache.scala 125:{53,53}]
  wire  _GEN_555 = 7'h20 == reqIndex ? way0Age_32 : _GEN_554; // @[DCache.scala 125:{53,53}]
  wire  _GEN_556 = 7'h21 == reqIndex ? way0Age_33 : _GEN_555; // @[DCache.scala 125:{53,53}]
  wire  _GEN_557 = 7'h22 == reqIndex ? way0Age_34 : _GEN_556; // @[DCache.scala 125:{53,53}]
  wire  _GEN_558 = 7'h23 == reqIndex ? way0Age_35 : _GEN_557; // @[DCache.scala 125:{53,53}]
  wire  _GEN_559 = 7'h24 == reqIndex ? way0Age_36 : _GEN_558; // @[DCache.scala 125:{53,53}]
  wire  _GEN_560 = 7'h25 == reqIndex ? way0Age_37 : _GEN_559; // @[DCache.scala 125:{53,53}]
  wire  _GEN_561 = 7'h26 == reqIndex ? way0Age_38 : _GEN_560; // @[DCache.scala 125:{53,53}]
  wire  _GEN_562 = 7'h27 == reqIndex ? way0Age_39 : _GEN_561; // @[DCache.scala 125:{53,53}]
  wire  _GEN_563 = 7'h28 == reqIndex ? way0Age_40 : _GEN_562; // @[DCache.scala 125:{53,53}]
  wire  _GEN_564 = 7'h29 == reqIndex ? way0Age_41 : _GEN_563; // @[DCache.scala 125:{53,53}]
  wire  _GEN_565 = 7'h2a == reqIndex ? way0Age_42 : _GEN_564; // @[DCache.scala 125:{53,53}]
  wire  _GEN_566 = 7'h2b == reqIndex ? way0Age_43 : _GEN_565; // @[DCache.scala 125:{53,53}]
  wire  _GEN_567 = 7'h2c == reqIndex ? way0Age_44 : _GEN_566; // @[DCache.scala 125:{53,53}]
  wire  _GEN_568 = 7'h2d == reqIndex ? way0Age_45 : _GEN_567; // @[DCache.scala 125:{53,53}]
  wire  _GEN_569 = 7'h2e == reqIndex ? way0Age_46 : _GEN_568; // @[DCache.scala 125:{53,53}]
  wire  _GEN_570 = 7'h2f == reqIndex ? way0Age_47 : _GEN_569; // @[DCache.scala 125:{53,53}]
  wire  _GEN_571 = 7'h30 == reqIndex ? way0Age_48 : _GEN_570; // @[DCache.scala 125:{53,53}]
  wire  _GEN_572 = 7'h31 == reqIndex ? way0Age_49 : _GEN_571; // @[DCache.scala 125:{53,53}]
  wire  _GEN_573 = 7'h32 == reqIndex ? way0Age_50 : _GEN_572; // @[DCache.scala 125:{53,53}]
  wire  _GEN_574 = 7'h33 == reqIndex ? way0Age_51 : _GEN_573; // @[DCache.scala 125:{53,53}]
  wire  _GEN_575 = 7'h34 == reqIndex ? way0Age_52 : _GEN_574; // @[DCache.scala 125:{53,53}]
  wire  _GEN_576 = 7'h35 == reqIndex ? way0Age_53 : _GEN_575; // @[DCache.scala 125:{53,53}]
  wire  _GEN_577 = 7'h36 == reqIndex ? way0Age_54 : _GEN_576; // @[DCache.scala 125:{53,53}]
  wire  _GEN_578 = 7'h37 == reqIndex ? way0Age_55 : _GEN_577; // @[DCache.scala 125:{53,53}]
  wire  _GEN_579 = 7'h38 == reqIndex ? way0Age_56 : _GEN_578; // @[DCache.scala 125:{53,53}]
  wire  _GEN_580 = 7'h39 == reqIndex ? way0Age_57 : _GEN_579; // @[DCache.scala 125:{53,53}]
  wire  _GEN_581 = 7'h3a == reqIndex ? way0Age_58 : _GEN_580; // @[DCache.scala 125:{53,53}]
  wire  _GEN_582 = 7'h3b == reqIndex ? way0Age_59 : _GEN_581; // @[DCache.scala 125:{53,53}]
  wire  _GEN_583 = 7'h3c == reqIndex ? way0Age_60 : _GEN_582; // @[DCache.scala 125:{53,53}]
  wire  _GEN_584 = 7'h3d == reqIndex ? way0Age_61 : _GEN_583; // @[DCache.scala 125:{53,53}]
  wire  _GEN_585 = 7'h3e == reqIndex ? way0Age_62 : _GEN_584; // @[DCache.scala 125:{53,53}]
  wire  _GEN_586 = 7'h3f == reqIndex ? way0Age_63 : _GEN_585; // @[DCache.scala 125:{53,53}]
  wire  _GEN_587 = 7'h40 == reqIndex ? way0Age_64 : _GEN_586; // @[DCache.scala 125:{53,53}]
  wire  _GEN_588 = 7'h41 == reqIndex ? way0Age_65 : _GEN_587; // @[DCache.scala 125:{53,53}]
  wire  _GEN_589 = 7'h42 == reqIndex ? way0Age_66 : _GEN_588; // @[DCache.scala 125:{53,53}]
  wire  _GEN_590 = 7'h43 == reqIndex ? way0Age_67 : _GEN_589; // @[DCache.scala 125:{53,53}]
  wire  _GEN_591 = 7'h44 == reqIndex ? way0Age_68 : _GEN_590; // @[DCache.scala 125:{53,53}]
  wire  _GEN_592 = 7'h45 == reqIndex ? way0Age_69 : _GEN_591; // @[DCache.scala 125:{53,53}]
  wire  _GEN_593 = 7'h46 == reqIndex ? way0Age_70 : _GEN_592; // @[DCache.scala 125:{53,53}]
  wire  _GEN_594 = 7'h47 == reqIndex ? way0Age_71 : _GEN_593; // @[DCache.scala 125:{53,53}]
  wire  _GEN_595 = 7'h48 == reqIndex ? way0Age_72 : _GEN_594; // @[DCache.scala 125:{53,53}]
  wire  _GEN_596 = 7'h49 == reqIndex ? way0Age_73 : _GEN_595; // @[DCache.scala 125:{53,53}]
  wire  _GEN_597 = 7'h4a == reqIndex ? way0Age_74 : _GEN_596; // @[DCache.scala 125:{53,53}]
  wire  _GEN_598 = 7'h4b == reqIndex ? way0Age_75 : _GEN_597; // @[DCache.scala 125:{53,53}]
  wire  _GEN_599 = 7'h4c == reqIndex ? way0Age_76 : _GEN_598; // @[DCache.scala 125:{53,53}]
  wire  _GEN_600 = 7'h4d == reqIndex ? way0Age_77 : _GEN_599; // @[DCache.scala 125:{53,53}]
  wire  _GEN_601 = 7'h4e == reqIndex ? way0Age_78 : _GEN_600; // @[DCache.scala 125:{53,53}]
  wire  _GEN_602 = 7'h4f == reqIndex ? way0Age_79 : _GEN_601; // @[DCache.scala 125:{53,53}]
  wire  _GEN_603 = 7'h50 == reqIndex ? way0Age_80 : _GEN_602; // @[DCache.scala 125:{53,53}]
  wire  _GEN_604 = 7'h51 == reqIndex ? way0Age_81 : _GEN_603; // @[DCache.scala 125:{53,53}]
  wire  _GEN_605 = 7'h52 == reqIndex ? way0Age_82 : _GEN_604; // @[DCache.scala 125:{53,53}]
  wire  _GEN_606 = 7'h53 == reqIndex ? way0Age_83 : _GEN_605; // @[DCache.scala 125:{53,53}]
  wire  _GEN_607 = 7'h54 == reqIndex ? way0Age_84 : _GEN_606; // @[DCache.scala 125:{53,53}]
  wire  _GEN_608 = 7'h55 == reqIndex ? way0Age_85 : _GEN_607; // @[DCache.scala 125:{53,53}]
  wire  _GEN_609 = 7'h56 == reqIndex ? way0Age_86 : _GEN_608; // @[DCache.scala 125:{53,53}]
  wire  _GEN_610 = 7'h57 == reqIndex ? way0Age_87 : _GEN_609; // @[DCache.scala 125:{53,53}]
  wire  _GEN_611 = 7'h58 == reqIndex ? way0Age_88 : _GEN_610; // @[DCache.scala 125:{53,53}]
  wire  _GEN_612 = 7'h59 == reqIndex ? way0Age_89 : _GEN_611; // @[DCache.scala 125:{53,53}]
  wire  _GEN_613 = 7'h5a == reqIndex ? way0Age_90 : _GEN_612; // @[DCache.scala 125:{53,53}]
  wire  _GEN_614 = 7'h5b == reqIndex ? way0Age_91 : _GEN_613; // @[DCache.scala 125:{53,53}]
  wire  _GEN_615 = 7'h5c == reqIndex ? way0Age_92 : _GEN_614; // @[DCache.scala 125:{53,53}]
  wire  _GEN_616 = 7'h5d == reqIndex ? way0Age_93 : _GEN_615; // @[DCache.scala 125:{53,53}]
  wire  _GEN_617 = 7'h5e == reqIndex ? way0Age_94 : _GEN_616; // @[DCache.scala 125:{53,53}]
  wire  _GEN_618 = 7'h5f == reqIndex ? way0Age_95 : _GEN_617; // @[DCache.scala 125:{53,53}]
  wire  _GEN_619 = 7'h60 == reqIndex ? way0Age_96 : _GEN_618; // @[DCache.scala 125:{53,53}]
  wire  _GEN_620 = 7'h61 == reqIndex ? way0Age_97 : _GEN_619; // @[DCache.scala 125:{53,53}]
  wire  _GEN_621 = 7'h62 == reqIndex ? way0Age_98 : _GEN_620; // @[DCache.scala 125:{53,53}]
  wire  _GEN_622 = 7'h63 == reqIndex ? way0Age_99 : _GEN_621; // @[DCache.scala 125:{53,53}]
  wire  _GEN_623 = 7'h64 == reqIndex ? way0Age_100 : _GEN_622; // @[DCache.scala 125:{53,53}]
  wire  _GEN_624 = 7'h65 == reqIndex ? way0Age_101 : _GEN_623; // @[DCache.scala 125:{53,53}]
  wire  _GEN_625 = 7'h66 == reqIndex ? way0Age_102 : _GEN_624; // @[DCache.scala 125:{53,53}]
  wire  _GEN_626 = 7'h67 == reqIndex ? way0Age_103 : _GEN_625; // @[DCache.scala 125:{53,53}]
  wire  _GEN_627 = 7'h68 == reqIndex ? way0Age_104 : _GEN_626; // @[DCache.scala 125:{53,53}]
  wire  _GEN_628 = 7'h69 == reqIndex ? way0Age_105 : _GEN_627; // @[DCache.scala 125:{53,53}]
  wire  _GEN_629 = 7'h6a == reqIndex ? way0Age_106 : _GEN_628; // @[DCache.scala 125:{53,53}]
  wire  _GEN_630 = 7'h6b == reqIndex ? way0Age_107 : _GEN_629; // @[DCache.scala 125:{53,53}]
  wire  _GEN_631 = 7'h6c == reqIndex ? way0Age_108 : _GEN_630; // @[DCache.scala 125:{53,53}]
  wire  _GEN_632 = 7'h6d == reqIndex ? way0Age_109 : _GEN_631; // @[DCache.scala 125:{53,53}]
  wire  _GEN_633 = 7'h6e == reqIndex ? way0Age_110 : _GEN_632; // @[DCache.scala 125:{53,53}]
  wire  _GEN_634 = 7'h6f == reqIndex ? way0Age_111 : _GEN_633; // @[DCache.scala 125:{53,53}]
  wire  _GEN_635 = 7'h70 == reqIndex ? way0Age_112 : _GEN_634; // @[DCache.scala 125:{53,53}]
  wire  _GEN_636 = 7'h71 == reqIndex ? way0Age_113 : _GEN_635; // @[DCache.scala 125:{53,53}]
  wire  _GEN_637 = 7'h72 == reqIndex ? way0Age_114 : _GEN_636; // @[DCache.scala 125:{53,53}]
  wire  _GEN_638 = 7'h73 == reqIndex ? way0Age_115 : _GEN_637; // @[DCache.scala 125:{53,53}]
  wire  _GEN_639 = 7'h74 == reqIndex ? way0Age_116 : _GEN_638; // @[DCache.scala 125:{53,53}]
  wire  _GEN_640 = 7'h75 == reqIndex ? way0Age_117 : _GEN_639; // @[DCache.scala 125:{53,53}]
  wire  _GEN_641 = 7'h76 == reqIndex ? way0Age_118 : _GEN_640; // @[DCache.scala 125:{53,53}]
  wire  _GEN_642 = 7'h77 == reqIndex ? way0Age_119 : _GEN_641; // @[DCache.scala 125:{53,53}]
  wire  _GEN_643 = 7'h78 == reqIndex ? way0Age_120 : _GEN_642; // @[DCache.scala 125:{53,53}]
  wire  _GEN_644 = 7'h79 == reqIndex ? way0Age_121 : _GEN_643; // @[DCache.scala 125:{53,53}]
  wire  _GEN_645 = 7'h7a == reqIndex ? way0Age_122 : _GEN_644; // @[DCache.scala 125:{53,53}]
  wire  _GEN_646 = 7'h7b == reqIndex ? way0Age_123 : _GEN_645; // @[DCache.scala 125:{53,53}]
  wire  _GEN_647 = 7'h7c == reqIndex ? way0Age_124 : _GEN_646; // @[DCache.scala 125:{53,53}]
  wire  _GEN_648 = 7'h7d == reqIndex ? way0Age_125 : _GEN_647; // @[DCache.scala 125:{53,53}]
  wire  _GEN_649 = 7'h7e == reqIndex ? way0Age_126 : _GEN_648; // @[DCache.scala 125:{53,53}]
  wire  _GEN_650 = 7'h7f == reqIndex ? way0Age_127 : _GEN_649; // @[DCache.scala 125:{53,53}]
  wire  ageWay0En = ~cacheHitEn & ~_GEN_650 & sHitEn; // @[DCache.scala 125:62]
  wire  cacheLineWay = ageWay0En ? 1'h0 : 1'h1; // @[DCache.scala 127:22]
  wire  _cacheDirtyEn_T = ~cacheLineWay; // @[DCache.scala 131:36]
  wire  sDirtyEn = state == 3'h2; // @[DCache.scala 130:24]
  wire  _GEN_780 = 7'h1 == reqIndex ? way0Dirty_1 : way0Dirty_0; // @[DCache.scala 131:{78,78}]
  wire  _GEN_781 = 7'h2 == reqIndex ? way0Dirty_2 : _GEN_780; // @[DCache.scala 131:{78,78}]
  wire  _GEN_782 = 7'h3 == reqIndex ? way0Dirty_3 : _GEN_781; // @[DCache.scala 131:{78,78}]
  wire  _GEN_783 = 7'h4 == reqIndex ? way0Dirty_4 : _GEN_782; // @[DCache.scala 131:{78,78}]
  wire  _GEN_784 = 7'h5 == reqIndex ? way0Dirty_5 : _GEN_783; // @[DCache.scala 131:{78,78}]
  wire  _GEN_785 = 7'h6 == reqIndex ? way0Dirty_6 : _GEN_784; // @[DCache.scala 131:{78,78}]
  wire  _GEN_786 = 7'h7 == reqIndex ? way0Dirty_7 : _GEN_785; // @[DCache.scala 131:{78,78}]
  wire  _GEN_787 = 7'h8 == reqIndex ? way0Dirty_8 : _GEN_786; // @[DCache.scala 131:{78,78}]
  wire  _GEN_788 = 7'h9 == reqIndex ? way0Dirty_9 : _GEN_787; // @[DCache.scala 131:{78,78}]
  wire  _GEN_789 = 7'ha == reqIndex ? way0Dirty_10 : _GEN_788; // @[DCache.scala 131:{78,78}]
  wire  _GEN_790 = 7'hb == reqIndex ? way0Dirty_11 : _GEN_789; // @[DCache.scala 131:{78,78}]
  wire  _GEN_791 = 7'hc == reqIndex ? way0Dirty_12 : _GEN_790; // @[DCache.scala 131:{78,78}]
  wire  _GEN_792 = 7'hd == reqIndex ? way0Dirty_13 : _GEN_791; // @[DCache.scala 131:{78,78}]
  wire  _GEN_793 = 7'he == reqIndex ? way0Dirty_14 : _GEN_792; // @[DCache.scala 131:{78,78}]
  wire  _GEN_794 = 7'hf == reqIndex ? way0Dirty_15 : _GEN_793; // @[DCache.scala 131:{78,78}]
  wire  _GEN_795 = 7'h10 == reqIndex ? way0Dirty_16 : _GEN_794; // @[DCache.scala 131:{78,78}]
  wire  _GEN_796 = 7'h11 == reqIndex ? way0Dirty_17 : _GEN_795; // @[DCache.scala 131:{78,78}]
  wire  _GEN_797 = 7'h12 == reqIndex ? way0Dirty_18 : _GEN_796; // @[DCache.scala 131:{78,78}]
  wire  _GEN_798 = 7'h13 == reqIndex ? way0Dirty_19 : _GEN_797; // @[DCache.scala 131:{78,78}]
  wire  _GEN_799 = 7'h14 == reqIndex ? way0Dirty_20 : _GEN_798; // @[DCache.scala 131:{78,78}]
  wire  _GEN_800 = 7'h15 == reqIndex ? way0Dirty_21 : _GEN_799; // @[DCache.scala 131:{78,78}]
  wire  _GEN_801 = 7'h16 == reqIndex ? way0Dirty_22 : _GEN_800; // @[DCache.scala 131:{78,78}]
  wire  _GEN_802 = 7'h17 == reqIndex ? way0Dirty_23 : _GEN_801; // @[DCache.scala 131:{78,78}]
  wire  _GEN_803 = 7'h18 == reqIndex ? way0Dirty_24 : _GEN_802; // @[DCache.scala 131:{78,78}]
  wire  _GEN_804 = 7'h19 == reqIndex ? way0Dirty_25 : _GEN_803; // @[DCache.scala 131:{78,78}]
  wire  _GEN_805 = 7'h1a == reqIndex ? way0Dirty_26 : _GEN_804; // @[DCache.scala 131:{78,78}]
  wire  _GEN_806 = 7'h1b == reqIndex ? way0Dirty_27 : _GEN_805; // @[DCache.scala 131:{78,78}]
  wire  _GEN_807 = 7'h1c == reqIndex ? way0Dirty_28 : _GEN_806; // @[DCache.scala 131:{78,78}]
  wire  _GEN_808 = 7'h1d == reqIndex ? way0Dirty_29 : _GEN_807; // @[DCache.scala 131:{78,78}]
  wire  _GEN_809 = 7'h1e == reqIndex ? way0Dirty_30 : _GEN_808; // @[DCache.scala 131:{78,78}]
  wire  _GEN_810 = 7'h1f == reqIndex ? way0Dirty_31 : _GEN_809; // @[DCache.scala 131:{78,78}]
  wire  _GEN_811 = 7'h20 == reqIndex ? way0Dirty_32 : _GEN_810; // @[DCache.scala 131:{78,78}]
  wire  _GEN_812 = 7'h21 == reqIndex ? way0Dirty_33 : _GEN_811; // @[DCache.scala 131:{78,78}]
  wire  _GEN_813 = 7'h22 == reqIndex ? way0Dirty_34 : _GEN_812; // @[DCache.scala 131:{78,78}]
  wire  _GEN_814 = 7'h23 == reqIndex ? way0Dirty_35 : _GEN_813; // @[DCache.scala 131:{78,78}]
  wire  _GEN_815 = 7'h24 == reqIndex ? way0Dirty_36 : _GEN_814; // @[DCache.scala 131:{78,78}]
  wire  _GEN_816 = 7'h25 == reqIndex ? way0Dirty_37 : _GEN_815; // @[DCache.scala 131:{78,78}]
  wire  _GEN_817 = 7'h26 == reqIndex ? way0Dirty_38 : _GEN_816; // @[DCache.scala 131:{78,78}]
  wire  _GEN_818 = 7'h27 == reqIndex ? way0Dirty_39 : _GEN_817; // @[DCache.scala 131:{78,78}]
  wire  _GEN_819 = 7'h28 == reqIndex ? way0Dirty_40 : _GEN_818; // @[DCache.scala 131:{78,78}]
  wire  _GEN_820 = 7'h29 == reqIndex ? way0Dirty_41 : _GEN_819; // @[DCache.scala 131:{78,78}]
  wire  _GEN_821 = 7'h2a == reqIndex ? way0Dirty_42 : _GEN_820; // @[DCache.scala 131:{78,78}]
  wire  _GEN_822 = 7'h2b == reqIndex ? way0Dirty_43 : _GEN_821; // @[DCache.scala 131:{78,78}]
  wire  _GEN_823 = 7'h2c == reqIndex ? way0Dirty_44 : _GEN_822; // @[DCache.scala 131:{78,78}]
  wire  _GEN_824 = 7'h2d == reqIndex ? way0Dirty_45 : _GEN_823; // @[DCache.scala 131:{78,78}]
  wire  _GEN_825 = 7'h2e == reqIndex ? way0Dirty_46 : _GEN_824; // @[DCache.scala 131:{78,78}]
  wire  _GEN_826 = 7'h2f == reqIndex ? way0Dirty_47 : _GEN_825; // @[DCache.scala 131:{78,78}]
  wire  _GEN_827 = 7'h30 == reqIndex ? way0Dirty_48 : _GEN_826; // @[DCache.scala 131:{78,78}]
  wire  _GEN_828 = 7'h31 == reqIndex ? way0Dirty_49 : _GEN_827; // @[DCache.scala 131:{78,78}]
  wire  _GEN_829 = 7'h32 == reqIndex ? way0Dirty_50 : _GEN_828; // @[DCache.scala 131:{78,78}]
  wire  _GEN_830 = 7'h33 == reqIndex ? way0Dirty_51 : _GEN_829; // @[DCache.scala 131:{78,78}]
  wire  _GEN_831 = 7'h34 == reqIndex ? way0Dirty_52 : _GEN_830; // @[DCache.scala 131:{78,78}]
  wire  _GEN_832 = 7'h35 == reqIndex ? way0Dirty_53 : _GEN_831; // @[DCache.scala 131:{78,78}]
  wire  _GEN_833 = 7'h36 == reqIndex ? way0Dirty_54 : _GEN_832; // @[DCache.scala 131:{78,78}]
  wire  _GEN_834 = 7'h37 == reqIndex ? way0Dirty_55 : _GEN_833; // @[DCache.scala 131:{78,78}]
  wire  _GEN_835 = 7'h38 == reqIndex ? way0Dirty_56 : _GEN_834; // @[DCache.scala 131:{78,78}]
  wire  _GEN_836 = 7'h39 == reqIndex ? way0Dirty_57 : _GEN_835; // @[DCache.scala 131:{78,78}]
  wire  _GEN_837 = 7'h3a == reqIndex ? way0Dirty_58 : _GEN_836; // @[DCache.scala 131:{78,78}]
  wire  _GEN_838 = 7'h3b == reqIndex ? way0Dirty_59 : _GEN_837; // @[DCache.scala 131:{78,78}]
  wire  _GEN_839 = 7'h3c == reqIndex ? way0Dirty_60 : _GEN_838; // @[DCache.scala 131:{78,78}]
  wire  _GEN_840 = 7'h3d == reqIndex ? way0Dirty_61 : _GEN_839; // @[DCache.scala 131:{78,78}]
  wire  _GEN_841 = 7'h3e == reqIndex ? way0Dirty_62 : _GEN_840; // @[DCache.scala 131:{78,78}]
  wire  _GEN_842 = 7'h3f == reqIndex ? way0Dirty_63 : _GEN_841; // @[DCache.scala 131:{78,78}]
  wire  _GEN_843 = 7'h40 == reqIndex ? way0Dirty_64 : _GEN_842; // @[DCache.scala 131:{78,78}]
  wire  _GEN_844 = 7'h41 == reqIndex ? way0Dirty_65 : _GEN_843; // @[DCache.scala 131:{78,78}]
  wire  _GEN_845 = 7'h42 == reqIndex ? way0Dirty_66 : _GEN_844; // @[DCache.scala 131:{78,78}]
  wire  _GEN_846 = 7'h43 == reqIndex ? way0Dirty_67 : _GEN_845; // @[DCache.scala 131:{78,78}]
  wire  _GEN_847 = 7'h44 == reqIndex ? way0Dirty_68 : _GEN_846; // @[DCache.scala 131:{78,78}]
  wire  _GEN_848 = 7'h45 == reqIndex ? way0Dirty_69 : _GEN_847; // @[DCache.scala 131:{78,78}]
  wire  _GEN_849 = 7'h46 == reqIndex ? way0Dirty_70 : _GEN_848; // @[DCache.scala 131:{78,78}]
  wire  _GEN_850 = 7'h47 == reqIndex ? way0Dirty_71 : _GEN_849; // @[DCache.scala 131:{78,78}]
  wire  _GEN_851 = 7'h48 == reqIndex ? way0Dirty_72 : _GEN_850; // @[DCache.scala 131:{78,78}]
  wire  _GEN_852 = 7'h49 == reqIndex ? way0Dirty_73 : _GEN_851; // @[DCache.scala 131:{78,78}]
  wire  _GEN_853 = 7'h4a == reqIndex ? way0Dirty_74 : _GEN_852; // @[DCache.scala 131:{78,78}]
  wire  _GEN_854 = 7'h4b == reqIndex ? way0Dirty_75 : _GEN_853; // @[DCache.scala 131:{78,78}]
  wire  _GEN_855 = 7'h4c == reqIndex ? way0Dirty_76 : _GEN_854; // @[DCache.scala 131:{78,78}]
  wire  _GEN_856 = 7'h4d == reqIndex ? way0Dirty_77 : _GEN_855; // @[DCache.scala 131:{78,78}]
  wire  _GEN_857 = 7'h4e == reqIndex ? way0Dirty_78 : _GEN_856; // @[DCache.scala 131:{78,78}]
  wire  _GEN_858 = 7'h4f == reqIndex ? way0Dirty_79 : _GEN_857; // @[DCache.scala 131:{78,78}]
  wire  _GEN_859 = 7'h50 == reqIndex ? way0Dirty_80 : _GEN_858; // @[DCache.scala 131:{78,78}]
  wire  _GEN_860 = 7'h51 == reqIndex ? way0Dirty_81 : _GEN_859; // @[DCache.scala 131:{78,78}]
  wire  _GEN_861 = 7'h52 == reqIndex ? way0Dirty_82 : _GEN_860; // @[DCache.scala 131:{78,78}]
  wire  _GEN_862 = 7'h53 == reqIndex ? way0Dirty_83 : _GEN_861; // @[DCache.scala 131:{78,78}]
  wire  _GEN_863 = 7'h54 == reqIndex ? way0Dirty_84 : _GEN_862; // @[DCache.scala 131:{78,78}]
  wire  _GEN_864 = 7'h55 == reqIndex ? way0Dirty_85 : _GEN_863; // @[DCache.scala 131:{78,78}]
  wire  _GEN_865 = 7'h56 == reqIndex ? way0Dirty_86 : _GEN_864; // @[DCache.scala 131:{78,78}]
  wire  _GEN_866 = 7'h57 == reqIndex ? way0Dirty_87 : _GEN_865; // @[DCache.scala 131:{78,78}]
  wire  _GEN_867 = 7'h58 == reqIndex ? way0Dirty_88 : _GEN_866; // @[DCache.scala 131:{78,78}]
  wire  _GEN_868 = 7'h59 == reqIndex ? way0Dirty_89 : _GEN_867; // @[DCache.scala 131:{78,78}]
  wire  _GEN_869 = 7'h5a == reqIndex ? way0Dirty_90 : _GEN_868; // @[DCache.scala 131:{78,78}]
  wire  _GEN_870 = 7'h5b == reqIndex ? way0Dirty_91 : _GEN_869; // @[DCache.scala 131:{78,78}]
  wire  _GEN_871 = 7'h5c == reqIndex ? way0Dirty_92 : _GEN_870; // @[DCache.scala 131:{78,78}]
  wire  _GEN_872 = 7'h5d == reqIndex ? way0Dirty_93 : _GEN_871; // @[DCache.scala 131:{78,78}]
  wire  _GEN_873 = 7'h5e == reqIndex ? way0Dirty_94 : _GEN_872; // @[DCache.scala 131:{78,78}]
  wire  _GEN_874 = 7'h5f == reqIndex ? way0Dirty_95 : _GEN_873; // @[DCache.scala 131:{78,78}]
  wire  _GEN_875 = 7'h60 == reqIndex ? way0Dirty_96 : _GEN_874; // @[DCache.scala 131:{78,78}]
  wire  _GEN_876 = 7'h61 == reqIndex ? way0Dirty_97 : _GEN_875; // @[DCache.scala 131:{78,78}]
  wire  _GEN_877 = 7'h62 == reqIndex ? way0Dirty_98 : _GEN_876; // @[DCache.scala 131:{78,78}]
  wire  _GEN_878 = 7'h63 == reqIndex ? way0Dirty_99 : _GEN_877; // @[DCache.scala 131:{78,78}]
  wire  _GEN_879 = 7'h64 == reqIndex ? way0Dirty_100 : _GEN_878; // @[DCache.scala 131:{78,78}]
  wire  _GEN_880 = 7'h65 == reqIndex ? way0Dirty_101 : _GEN_879; // @[DCache.scala 131:{78,78}]
  wire  _GEN_881 = 7'h66 == reqIndex ? way0Dirty_102 : _GEN_880; // @[DCache.scala 131:{78,78}]
  wire  _GEN_882 = 7'h67 == reqIndex ? way0Dirty_103 : _GEN_881; // @[DCache.scala 131:{78,78}]
  wire  _GEN_883 = 7'h68 == reqIndex ? way0Dirty_104 : _GEN_882; // @[DCache.scala 131:{78,78}]
  wire  _GEN_884 = 7'h69 == reqIndex ? way0Dirty_105 : _GEN_883; // @[DCache.scala 131:{78,78}]
  wire  _GEN_885 = 7'h6a == reqIndex ? way0Dirty_106 : _GEN_884; // @[DCache.scala 131:{78,78}]
  wire  _GEN_886 = 7'h6b == reqIndex ? way0Dirty_107 : _GEN_885; // @[DCache.scala 131:{78,78}]
  wire  _GEN_887 = 7'h6c == reqIndex ? way0Dirty_108 : _GEN_886; // @[DCache.scala 131:{78,78}]
  wire  _GEN_888 = 7'h6d == reqIndex ? way0Dirty_109 : _GEN_887; // @[DCache.scala 131:{78,78}]
  wire  _GEN_889 = 7'h6e == reqIndex ? way0Dirty_110 : _GEN_888; // @[DCache.scala 131:{78,78}]
  wire  _GEN_890 = 7'h6f == reqIndex ? way0Dirty_111 : _GEN_889; // @[DCache.scala 131:{78,78}]
  wire  _GEN_891 = 7'h70 == reqIndex ? way0Dirty_112 : _GEN_890; // @[DCache.scala 131:{78,78}]
  wire  _GEN_892 = 7'h71 == reqIndex ? way0Dirty_113 : _GEN_891; // @[DCache.scala 131:{78,78}]
  wire  _GEN_893 = 7'h72 == reqIndex ? way0Dirty_114 : _GEN_892; // @[DCache.scala 131:{78,78}]
  wire  _GEN_894 = 7'h73 == reqIndex ? way0Dirty_115 : _GEN_893; // @[DCache.scala 131:{78,78}]
  wire  _GEN_895 = 7'h74 == reqIndex ? way0Dirty_116 : _GEN_894; // @[DCache.scala 131:{78,78}]
  wire  _GEN_896 = 7'h75 == reqIndex ? way0Dirty_117 : _GEN_895; // @[DCache.scala 131:{78,78}]
  wire  _GEN_897 = 7'h76 == reqIndex ? way0Dirty_118 : _GEN_896; // @[DCache.scala 131:{78,78}]
  wire  _GEN_898 = 7'h77 == reqIndex ? way0Dirty_119 : _GEN_897; // @[DCache.scala 131:{78,78}]
  wire  _GEN_899 = 7'h78 == reqIndex ? way0Dirty_120 : _GEN_898; // @[DCache.scala 131:{78,78}]
  wire  _GEN_900 = 7'h79 == reqIndex ? way0Dirty_121 : _GEN_899; // @[DCache.scala 131:{78,78}]
  wire  _GEN_901 = 7'h7a == reqIndex ? way0Dirty_122 : _GEN_900; // @[DCache.scala 131:{78,78}]
  wire  _GEN_902 = 7'h7b == reqIndex ? way0Dirty_123 : _GEN_901; // @[DCache.scala 131:{78,78}]
  wire  _GEN_903 = 7'h7c == reqIndex ? way0Dirty_124 : _GEN_902; // @[DCache.scala 131:{78,78}]
  wire  _GEN_904 = 7'h7d == reqIndex ? way0Dirty_125 : _GEN_903; // @[DCache.scala 131:{78,78}]
  wire  _GEN_905 = 7'h7e == reqIndex ? way0Dirty_126 : _GEN_904; // @[DCache.scala 131:{78,78}]
  wire  _GEN_906 = 7'h7f == reqIndex ? way0Dirty_127 : _GEN_905; // @[DCache.scala 131:{78,78}]
  wire  _GEN_908 = 7'h1 == reqIndex ? way1Dirty_1 : way1Dirty_0; // @[DCache.scala 132:{54,54}]
  wire  _GEN_909 = 7'h2 == reqIndex ? way1Dirty_2 : _GEN_908; // @[DCache.scala 132:{54,54}]
  wire  _GEN_910 = 7'h3 == reqIndex ? way1Dirty_3 : _GEN_909; // @[DCache.scala 132:{54,54}]
  wire  _GEN_911 = 7'h4 == reqIndex ? way1Dirty_4 : _GEN_910; // @[DCache.scala 132:{54,54}]
  wire  _GEN_912 = 7'h5 == reqIndex ? way1Dirty_5 : _GEN_911; // @[DCache.scala 132:{54,54}]
  wire  _GEN_913 = 7'h6 == reqIndex ? way1Dirty_6 : _GEN_912; // @[DCache.scala 132:{54,54}]
  wire  _GEN_914 = 7'h7 == reqIndex ? way1Dirty_7 : _GEN_913; // @[DCache.scala 132:{54,54}]
  wire  _GEN_915 = 7'h8 == reqIndex ? way1Dirty_8 : _GEN_914; // @[DCache.scala 132:{54,54}]
  wire  _GEN_916 = 7'h9 == reqIndex ? way1Dirty_9 : _GEN_915; // @[DCache.scala 132:{54,54}]
  wire  _GEN_917 = 7'ha == reqIndex ? way1Dirty_10 : _GEN_916; // @[DCache.scala 132:{54,54}]
  wire  _GEN_918 = 7'hb == reqIndex ? way1Dirty_11 : _GEN_917; // @[DCache.scala 132:{54,54}]
  wire  _GEN_919 = 7'hc == reqIndex ? way1Dirty_12 : _GEN_918; // @[DCache.scala 132:{54,54}]
  wire  _GEN_920 = 7'hd == reqIndex ? way1Dirty_13 : _GEN_919; // @[DCache.scala 132:{54,54}]
  wire  _GEN_921 = 7'he == reqIndex ? way1Dirty_14 : _GEN_920; // @[DCache.scala 132:{54,54}]
  wire  _GEN_922 = 7'hf == reqIndex ? way1Dirty_15 : _GEN_921; // @[DCache.scala 132:{54,54}]
  wire  _GEN_923 = 7'h10 == reqIndex ? way1Dirty_16 : _GEN_922; // @[DCache.scala 132:{54,54}]
  wire  _GEN_924 = 7'h11 == reqIndex ? way1Dirty_17 : _GEN_923; // @[DCache.scala 132:{54,54}]
  wire  _GEN_925 = 7'h12 == reqIndex ? way1Dirty_18 : _GEN_924; // @[DCache.scala 132:{54,54}]
  wire  _GEN_926 = 7'h13 == reqIndex ? way1Dirty_19 : _GEN_925; // @[DCache.scala 132:{54,54}]
  wire  _GEN_927 = 7'h14 == reqIndex ? way1Dirty_20 : _GEN_926; // @[DCache.scala 132:{54,54}]
  wire  _GEN_928 = 7'h15 == reqIndex ? way1Dirty_21 : _GEN_927; // @[DCache.scala 132:{54,54}]
  wire  _GEN_929 = 7'h16 == reqIndex ? way1Dirty_22 : _GEN_928; // @[DCache.scala 132:{54,54}]
  wire  _GEN_930 = 7'h17 == reqIndex ? way1Dirty_23 : _GEN_929; // @[DCache.scala 132:{54,54}]
  wire  _GEN_931 = 7'h18 == reqIndex ? way1Dirty_24 : _GEN_930; // @[DCache.scala 132:{54,54}]
  wire  _GEN_932 = 7'h19 == reqIndex ? way1Dirty_25 : _GEN_931; // @[DCache.scala 132:{54,54}]
  wire  _GEN_933 = 7'h1a == reqIndex ? way1Dirty_26 : _GEN_932; // @[DCache.scala 132:{54,54}]
  wire  _GEN_934 = 7'h1b == reqIndex ? way1Dirty_27 : _GEN_933; // @[DCache.scala 132:{54,54}]
  wire  _GEN_935 = 7'h1c == reqIndex ? way1Dirty_28 : _GEN_934; // @[DCache.scala 132:{54,54}]
  wire  _GEN_936 = 7'h1d == reqIndex ? way1Dirty_29 : _GEN_935; // @[DCache.scala 132:{54,54}]
  wire  _GEN_937 = 7'h1e == reqIndex ? way1Dirty_30 : _GEN_936; // @[DCache.scala 132:{54,54}]
  wire  _GEN_938 = 7'h1f == reqIndex ? way1Dirty_31 : _GEN_937; // @[DCache.scala 132:{54,54}]
  wire  _GEN_939 = 7'h20 == reqIndex ? way1Dirty_32 : _GEN_938; // @[DCache.scala 132:{54,54}]
  wire  _GEN_940 = 7'h21 == reqIndex ? way1Dirty_33 : _GEN_939; // @[DCache.scala 132:{54,54}]
  wire  _GEN_941 = 7'h22 == reqIndex ? way1Dirty_34 : _GEN_940; // @[DCache.scala 132:{54,54}]
  wire  _GEN_942 = 7'h23 == reqIndex ? way1Dirty_35 : _GEN_941; // @[DCache.scala 132:{54,54}]
  wire  _GEN_943 = 7'h24 == reqIndex ? way1Dirty_36 : _GEN_942; // @[DCache.scala 132:{54,54}]
  wire  _GEN_944 = 7'h25 == reqIndex ? way1Dirty_37 : _GEN_943; // @[DCache.scala 132:{54,54}]
  wire  _GEN_945 = 7'h26 == reqIndex ? way1Dirty_38 : _GEN_944; // @[DCache.scala 132:{54,54}]
  wire  _GEN_946 = 7'h27 == reqIndex ? way1Dirty_39 : _GEN_945; // @[DCache.scala 132:{54,54}]
  wire  _GEN_947 = 7'h28 == reqIndex ? way1Dirty_40 : _GEN_946; // @[DCache.scala 132:{54,54}]
  wire  _GEN_948 = 7'h29 == reqIndex ? way1Dirty_41 : _GEN_947; // @[DCache.scala 132:{54,54}]
  wire  _GEN_949 = 7'h2a == reqIndex ? way1Dirty_42 : _GEN_948; // @[DCache.scala 132:{54,54}]
  wire  _GEN_950 = 7'h2b == reqIndex ? way1Dirty_43 : _GEN_949; // @[DCache.scala 132:{54,54}]
  wire  _GEN_951 = 7'h2c == reqIndex ? way1Dirty_44 : _GEN_950; // @[DCache.scala 132:{54,54}]
  wire  _GEN_952 = 7'h2d == reqIndex ? way1Dirty_45 : _GEN_951; // @[DCache.scala 132:{54,54}]
  wire  _GEN_953 = 7'h2e == reqIndex ? way1Dirty_46 : _GEN_952; // @[DCache.scala 132:{54,54}]
  wire  _GEN_954 = 7'h2f == reqIndex ? way1Dirty_47 : _GEN_953; // @[DCache.scala 132:{54,54}]
  wire  _GEN_955 = 7'h30 == reqIndex ? way1Dirty_48 : _GEN_954; // @[DCache.scala 132:{54,54}]
  wire  _GEN_956 = 7'h31 == reqIndex ? way1Dirty_49 : _GEN_955; // @[DCache.scala 132:{54,54}]
  wire  _GEN_957 = 7'h32 == reqIndex ? way1Dirty_50 : _GEN_956; // @[DCache.scala 132:{54,54}]
  wire  _GEN_958 = 7'h33 == reqIndex ? way1Dirty_51 : _GEN_957; // @[DCache.scala 132:{54,54}]
  wire  _GEN_959 = 7'h34 == reqIndex ? way1Dirty_52 : _GEN_958; // @[DCache.scala 132:{54,54}]
  wire  _GEN_960 = 7'h35 == reqIndex ? way1Dirty_53 : _GEN_959; // @[DCache.scala 132:{54,54}]
  wire  _GEN_961 = 7'h36 == reqIndex ? way1Dirty_54 : _GEN_960; // @[DCache.scala 132:{54,54}]
  wire  _GEN_962 = 7'h37 == reqIndex ? way1Dirty_55 : _GEN_961; // @[DCache.scala 132:{54,54}]
  wire  _GEN_963 = 7'h38 == reqIndex ? way1Dirty_56 : _GEN_962; // @[DCache.scala 132:{54,54}]
  wire  _GEN_964 = 7'h39 == reqIndex ? way1Dirty_57 : _GEN_963; // @[DCache.scala 132:{54,54}]
  wire  _GEN_965 = 7'h3a == reqIndex ? way1Dirty_58 : _GEN_964; // @[DCache.scala 132:{54,54}]
  wire  _GEN_966 = 7'h3b == reqIndex ? way1Dirty_59 : _GEN_965; // @[DCache.scala 132:{54,54}]
  wire  _GEN_967 = 7'h3c == reqIndex ? way1Dirty_60 : _GEN_966; // @[DCache.scala 132:{54,54}]
  wire  _GEN_968 = 7'h3d == reqIndex ? way1Dirty_61 : _GEN_967; // @[DCache.scala 132:{54,54}]
  wire  _GEN_969 = 7'h3e == reqIndex ? way1Dirty_62 : _GEN_968; // @[DCache.scala 132:{54,54}]
  wire  _GEN_970 = 7'h3f == reqIndex ? way1Dirty_63 : _GEN_969; // @[DCache.scala 132:{54,54}]
  wire  _GEN_971 = 7'h40 == reqIndex ? way1Dirty_64 : _GEN_970; // @[DCache.scala 132:{54,54}]
  wire  _GEN_972 = 7'h41 == reqIndex ? way1Dirty_65 : _GEN_971; // @[DCache.scala 132:{54,54}]
  wire  _GEN_973 = 7'h42 == reqIndex ? way1Dirty_66 : _GEN_972; // @[DCache.scala 132:{54,54}]
  wire  _GEN_974 = 7'h43 == reqIndex ? way1Dirty_67 : _GEN_973; // @[DCache.scala 132:{54,54}]
  wire  _GEN_975 = 7'h44 == reqIndex ? way1Dirty_68 : _GEN_974; // @[DCache.scala 132:{54,54}]
  wire  _GEN_976 = 7'h45 == reqIndex ? way1Dirty_69 : _GEN_975; // @[DCache.scala 132:{54,54}]
  wire  _GEN_977 = 7'h46 == reqIndex ? way1Dirty_70 : _GEN_976; // @[DCache.scala 132:{54,54}]
  wire  _GEN_978 = 7'h47 == reqIndex ? way1Dirty_71 : _GEN_977; // @[DCache.scala 132:{54,54}]
  wire  _GEN_979 = 7'h48 == reqIndex ? way1Dirty_72 : _GEN_978; // @[DCache.scala 132:{54,54}]
  wire  _GEN_980 = 7'h49 == reqIndex ? way1Dirty_73 : _GEN_979; // @[DCache.scala 132:{54,54}]
  wire  _GEN_981 = 7'h4a == reqIndex ? way1Dirty_74 : _GEN_980; // @[DCache.scala 132:{54,54}]
  wire  _GEN_982 = 7'h4b == reqIndex ? way1Dirty_75 : _GEN_981; // @[DCache.scala 132:{54,54}]
  wire  _GEN_983 = 7'h4c == reqIndex ? way1Dirty_76 : _GEN_982; // @[DCache.scala 132:{54,54}]
  wire  _GEN_984 = 7'h4d == reqIndex ? way1Dirty_77 : _GEN_983; // @[DCache.scala 132:{54,54}]
  wire  _GEN_985 = 7'h4e == reqIndex ? way1Dirty_78 : _GEN_984; // @[DCache.scala 132:{54,54}]
  wire  _GEN_986 = 7'h4f == reqIndex ? way1Dirty_79 : _GEN_985; // @[DCache.scala 132:{54,54}]
  wire  _GEN_987 = 7'h50 == reqIndex ? way1Dirty_80 : _GEN_986; // @[DCache.scala 132:{54,54}]
  wire  _GEN_988 = 7'h51 == reqIndex ? way1Dirty_81 : _GEN_987; // @[DCache.scala 132:{54,54}]
  wire  _GEN_989 = 7'h52 == reqIndex ? way1Dirty_82 : _GEN_988; // @[DCache.scala 132:{54,54}]
  wire  _GEN_990 = 7'h53 == reqIndex ? way1Dirty_83 : _GEN_989; // @[DCache.scala 132:{54,54}]
  wire  _GEN_991 = 7'h54 == reqIndex ? way1Dirty_84 : _GEN_990; // @[DCache.scala 132:{54,54}]
  wire  _GEN_992 = 7'h55 == reqIndex ? way1Dirty_85 : _GEN_991; // @[DCache.scala 132:{54,54}]
  wire  _GEN_993 = 7'h56 == reqIndex ? way1Dirty_86 : _GEN_992; // @[DCache.scala 132:{54,54}]
  wire  _GEN_994 = 7'h57 == reqIndex ? way1Dirty_87 : _GEN_993; // @[DCache.scala 132:{54,54}]
  wire  _GEN_995 = 7'h58 == reqIndex ? way1Dirty_88 : _GEN_994; // @[DCache.scala 132:{54,54}]
  wire  _GEN_996 = 7'h59 == reqIndex ? way1Dirty_89 : _GEN_995; // @[DCache.scala 132:{54,54}]
  wire  _GEN_997 = 7'h5a == reqIndex ? way1Dirty_90 : _GEN_996; // @[DCache.scala 132:{54,54}]
  wire  _GEN_998 = 7'h5b == reqIndex ? way1Dirty_91 : _GEN_997; // @[DCache.scala 132:{54,54}]
  wire  _GEN_999 = 7'h5c == reqIndex ? way1Dirty_92 : _GEN_998; // @[DCache.scala 132:{54,54}]
  wire  _GEN_1000 = 7'h5d == reqIndex ? way1Dirty_93 : _GEN_999; // @[DCache.scala 132:{54,54}]
  wire  _GEN_1001 = 7'h5e == reqIndex ? way1Dirty_94 : _GEN_1000; // @[DCache.scala 132:{54,54}]
  wire  _GEN_1002 = 7'h5f == reqIndex ? way1Dirty_95 : _GEN_1001; // @[DCache.scala 132:{54,54}]
  wire  _GEN_1003 = 7'h60 == reqIndex ? way1Dirty_96 : _GEN_1002; // @[DCache.scala 132:{54,54}]
  wire  _GEN_1004 = 7'h61 == reqIndex ? way1Dirty_97 : _GEN_1003; // @[DCache.scala 132:{54,54}]
  wire  _GEN_1005 = 7'h62 == reqIndex ? way1Dirty_98 : _GEN_1004; // @[DCache.scala 132:{54,54}]
  wire  _GEN_1006 = 7'h63 == reqIndex ? way1Dirty_99 : _GEN_1005; // @[DCache.scala 132:{54,54}]
  wire  _GEN_1007 = 7'h64 == reqIndex ? way1Dirty_100 : _GEN_1006; // @[DCache.scala 132:{54,54}]
  wire  _GEN_1008 = 7'h65 == reqIndex ? way1Dirty_101 : _GEN_1007; // @[DCache.scala 132:{54,54}]
  wire  _GEN_1009 = 7'h66 == reqIndex ? way1Dirty_102 : _GEN_1008; // @[DCache.scala 132:{54,54}]
  wire  _GEN_1010 = 7'h67 == reqIndex ? way1Dirty_103 : _GEN_1009; // @[DCache.scala 132:{54,54}]
  wire  _GEN_1011 = 7'h68 == reqIndex ? way1Dirty_104 : _GEN_1010; // @[DCache.scala 132:{54,54}]
  wire  _GEN_1012 = 7'h69 == reqIndex ? way1Dirty_105 : _GEN_1011; // @[DCache.scala 132:{54,54}]
  wire  _GEN_1013 = 7'h6a == reqIndex ? way1Dirty_106 : _GEN_1012; // @[DCache.scala 132:{54,54}]
  wire  _GEN_1014 = 7'h6b == reqIndex ? way1Dirty_107 : _GEN_1013; // @[DCache.scala 132:{54,54}]
  wire  _GEN_1015 = 7'h6c == reqIndex ? way1Dirty_108 : _GEN_1014; // @[DCache.scala 132:{54,54}]
  wire  _GEN_1016 = 7'h6d == reqIndex ? way1Dirty_109 : _GEN_1015; // @[DCache.scala 132:{54,54}]
  wire  _GEN_1017 = 7'h6e == reqIndex ? way1Dirty_110 : _GEN_1016; // @[DCache.scala 132:{54,54}]
  wire  _GEN_1018 = 7'h6f == reqIndex ? way1Dirty_111 : _GEN_1017; // @[DCache.scala 132:{54,54}]
  wire  _GEN_1019 = 7'h70 == reqIndex ? way1Dirty_112 : _GEN_1018; // @[DCache.scala 132:{54,54}]
  wire  _GEN_1020 = 7'h71 == reqIndex ? way1Dirty_113 : _GEN_1019; // @[DCache.scala 132:{54,54}]
  wire  _GEN_1021 = 7'h72 == reqIndex ? way1Dirty_114 : _GEN_1020; // @[DCache.scala 132:{54,54}]
  wire  _GEN_1022 = 7'h73 == reqIndex ? way1Dirty_115 : _GEN_1021; // @[DCache.scala 132:{54,54}]
  wire  _GEN_1023 = 7'h74 == reqIndex ? way1Dirty_116 : _GEN_1022; // @[DCache.scala 132:{54,54}]
  wire  _GEN_1024 = 7'h75 == reqIndex ? way1Dirty_117 : _GEN_1023; // @[DCache.scala 132:{54,54}]
  wire  _GEN_1025 = 7'h76 == reqIndex ? way1Dirty_118 : _GEN_1024; // @[DCache.scala 132:{54,54}]
  wire  _GEN_1026 = 7'h77 == reqIndex ? way1Dirty_119 : _GEN_1025; // @[DCache.scala 132:{54,54}]
  wire  _GEN_1027 = 7'h78 == reqIndex ? way1Dirty_120 : _GEN_1026; // @[DCache.scala 132:{54,54}]
  wire  _GEN_1028 = 7'h79 == reqIndex ? way1Dirty_121 : _GEN_1027; // @[DCache.scala 132:{54,54}]
  wire  _GEN_1029 = 7'h7a == reqIndex ? way1Dirty_122 : _GEN_1028; // @[DCache.scala 132:{54,54}]
  wire  _GEN_1030 = 7'h7b == reqIndex ? way1Dirty_123 : _GEN_1029; // @[DCache.scala 132:{54,54}]
  wire  _GEN_1031 = 7'h7c == reqIndex ? way1Dirty_124 : _GEN_1030; // @[DCache.scala 132:{54,54}]
  wire  _GEN_1032 = 7'h7d == reqIndex ? way1Dirty_125 : _GEN_1031; // @[DCache.scala 132:{54,54}]
  wire  _GEN_1033 = 7'h7e == reqIndex ? way1Dirty_126 : _GEN_1032; // @[DCache.scala 132:{54,54}]
  wire  _GEN_1034 = 7'h7f == reqIndex ? way1Dirty_127 : _GEN_1033; // @[DCache.scala 132:{54,54}]
  wire  _cacheDirtyEn_T_4 = sDirtyEn & _GEN_1034; // @[DCache.scala 132:30]
  wire  cacheDirtyEn = ~cacheLineWay ? sDirtyEn & _GEN_906 : _cacheDirtyEn_T_4; // @[DCache.scala 131:22]
  wire [2:0] _GEN_2 = cacheDirtyEn ? 3'h3 : 3'h4; // @[DCache.scala 95:28 96:15 98:15]
  wire [2:0] _GEN_3 = io_out_data_ready ? 3'h4 : state; // @[DCache.scala 102:30 103:15 46:22]
  wire  sCacheWEn = state == 3'h4; // @[DCache.scala 135:26]
  reg  cacheWriteEn_REG; // @[DCache.scala 164:41]
  wire  cacheWriteEn = sCacheWEn & cacheWriteEn_REG; // @[DCache.scala 164:22]
  wire [2:0] _GEN_4 = cacheWriteEn ? 3'h5 : state; // @[DCache.scala 107:28 108:15 46:22]
  wire [2:0] _GEN_5 = 3'h5 == state ? 3'h0 : state; // @[DCache.scala 112:13 81:17 46:22]
  wire [2:0] _GEN_6 = 3'h4 == state ? _GEN_4 : _GEN_5; // @[DCache.scala 81:17]
  wire [2:0] _GEN_7 = 3'h3 == state ? _GEN_3 : _GEN_6; // @[DCache.scala 81:17]
  wire [7:0] _cacheIndex_T_1 = {1'h0,reqIndex}; // @[Cat.scala 31:58]
  wire [7:0] _cacheIndex_T_2 = {1'h1,reqIndex}; // @[Cat.scala 31:58]
  wire [7:0] _cacheIndex_T_3 = _cacheDirtyEn_T ? _cacheIndex_T_1 : _cacheIndex_T_2; // @[DCache.scala 128:20]
  wire  sWriteEn = state == 3'h3; // @[DCache.scala 134:24]
  wire [127:0] cacheRData = req_Q;
  wire [127:0] cacheWData = cacheHitEn ? cacheRData : io_out_data_read; // @[DCache.scala 166:23]
  wire [191:0] _wData_T_2 = {io_dmem_data_write,cacheWData[63:0]}; // @[Cat.scala 31:58]
  wire [191:0] _wData_T_4 = {cacheWData[127:64],io_dmem_data_write}; // @[Cat.scala 31:58]
  wire [191:0] wData = reqOff[3] ? _wData_T_2 : _wData_T_4; // @[DCache.scala 167:18]
  wire [191:0] _valid_WData_T = io_dmem_data_req ? wData : {{64'd0}, io_out_data_read}; // @[DCache.scala 169:21]
  wire  sDoneEn = state == 3'h5; // @[DCache.scala 172:23]
  wire  _GEN_3595 = 7'h0 == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1291 = 7'h0 == reqIndex | way0V_0; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3596 = 7'h1 == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1292 = 7'h1 == reqIndex | way0V_1; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3597 = 7'h2 == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1293 = 7'h2 == reqIndex | way0V_2; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3598 = 7'h3 == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1294 = 7'h3 == reqIndex | way0V_3; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3599 = 7'h4 == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1295 = 7'h4 == reqIndex | way0V_4; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3600 = 7'h5 == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1296 = 7'h5 == reqIndex | way0V_5; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3601 = 7'h6 == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1297 = 7'h6 == reqIndex | way0V_6; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3602 = 7'h7 == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1298 = 7'h7 == reqIndex | way0V_7; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3603 = 7'h8 == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1299 = 7'h8 == reqIndex | way0V_8; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3604 = 7'h9 == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1300 = 7'h9 == reqIndex | way0V_9; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3605 = 7'ha == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1301 = 7'ha == reqIndex | way0V_10; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3606 = 7'hb == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1302 = 7'hb == reqIndex | way0V_11; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3607 = 7'hc == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1303 = 7'hc == reqIndex | way0V_12; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3608 = 7'hd == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1304 = 7'hd == reqIndex | way0V_13; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3609 = 7'he == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1305 = 7'he == reqIndex | way0V_14; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3610 = 7'hf == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1306 = 7'hf == reqIndex | way0V_15; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3611 = 7'h10 == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1307 = 7'h10 == reqIndex | way0V_16; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3612 = 7'h11 == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1308 = 7'h11 == reqIndex | way0V_17; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3613 = 7'h12 == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1309 = 7'h12 == reqIndex | way0V_18; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3614 = 7'h13 == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1310 = 7'h13 == reqIndex | way0V_19; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3615 = 7'h14 == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1311 = 7'h14 == reqIndex | way0V_20; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3616 = 7'h15 == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1312 = 7'h15 == reqIndex | way0V_21; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3617 = 7'h16 == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1313 = 7'h16 == reqIndex | way0V_22; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3618 = 7'h17 == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1314 = 7'h17 == reqIndex | way0V_23; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3619 = 7'h18 == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1315 = 7'h18 == reqIndex | way0V_24; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3620 = 7'h19 == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1316 = 7'h19 == reqIndex | way0V_25; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3621 = 7'h1a == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1317 = 7'h1a == reqIndex | way0V_26; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3622 = 7'h1b == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1318 = 7'h1b == reqIndex | way0V_27; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3623 = 7'h1c == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1319 = 7'h1c == reqIndex | way0V_28; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3624 = 7'h1d == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1320 = 7'h1d == reqIndex | way0V_29; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3625 = 7'h1e == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1321 = 7'h1e == reqIndex | way0V_30; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3626 = 7'h1f == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1322 = 7'h1f == reqIndex | way0V_31; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3627 = 7'h20 == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1323 = 7'h20 == reqIndex | way0V_32; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3628 = 7'h21 == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1324 = 7'h21 == reqIndex | way0V_33; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3629 = 7'h22 == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1325 = 7'h22 == reqIndex | way0V_34; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3630 = 7'h23 == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1326 = 7'h23 == reqIndex | way0V_35; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3631 = 7'h24 == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1327 = 7'h24 == reqIndex | way0V_36; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3632 = 7'h25 == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1328 = 7'h25 == reqIndex | way0V_37; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3633 = 7'h26 == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1329 = 7'h26 == reqIndex | way0V_38; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3634 = 7'h27 == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1330 = 7'h27 == reqIndex | way0V_39; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3635 = 7'h28 == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1331 = 7'h28 == reqIndex | way0V_40; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3636 = 7'h29 == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1332 = 7'h29 == reqIndex | way0V_41; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3637 = 7'h2a == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1333 = 7'h2a == reqIndex | way0V_42; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3638 = 7'h2b == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1334 = 7'h2b == reqIndex | way0V_43; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3639 = 7'h2c == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1335 = 7'h2c == reqIndex | way0V_44; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3640 = 7'h2d == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1336 = 7'h2d == reqIndex | way0V_45; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3641 = 7'h2e == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1337 = 7'h2e == reqIndex | way0V_46; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3642 = 7'h2f == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1338 = 7'h2f == reqIndex | way0V_47; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3643 = 7'h30 == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1339 = 7'h30 == reqIndex | way0V_48; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3644 = 7'h31 == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1340 = 7'h31 == reqIndex | way0V_49; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3645 = 7'h32 == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1341 = 7'h32 == reqIndex | way0V_50; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3646 = 7'h33 == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1342 = 7'h33 == reqIndex | way0V_51; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3647 = 7'h34 == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1343 = 7'h34 == reqIndex | way0V_52; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3648 = 7'h35 == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1344 = 7'h35 == reqIndex | way0V_53; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3649 = 7'h36 == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1345 = 7'h36 == reqIndex | way0V_54; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3650 = 7'h37 == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1346 = 7'h37 == reqIndex | way0V_55; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3651 = 7'h38 == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1347 = 7'h38 == reqIndex | way0V_56; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3652 = 7'h39 == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1348 = 7'h39 == reqIndex | way0V_57; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3653 = 7'h3a == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1349 = 7'h3a == reqIndex | way0V_58; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3654 = 7'h3b == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1350 = 7'h3b == reqIndex | way0V_59; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3655 = 7'h3c == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1351 = 7'h3c == reqIndex | way0V_60; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3656 = 7'h3d == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1352 = 7'h3d == reqIndex | way0V_61; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3657 = 7'h3e == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1353 = 7'h3e == reqIndex | way0V_62; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3658 = 7'h3f == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1354 = 7'h3f == reqIndex | way0V_63; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3659 = 7'h40 == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1355 = 7'h40 == reqIndex | way0V_64; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3660 = 7'h41 == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1356 = 7'h41 == reqIndex | way0V_65; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3661 = 7'h42 == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1357 = 7'h42 == reqIndex | way0V_66; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3662 = 7'h43 == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1358 = 7'h43 == reqIndex | way0V_67; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3663 = 7'h44 == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1359 = 7'h44 == reqIndex | way0V_68; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3664 = 7'h45 == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1360 = 7'h45 == reqIndex | way0V_69; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3665 = 7'h46 == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1361 = 7'h46 == reqIndex | way0V_70; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3666 = 7'h47 == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1362 = 7'h47 == reqIndex | way0V_71; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3667 = 7'h48 == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1363 = 7'h48 == reqIndex | way0V_72; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3668 = 7'h49 == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1364 = 7'h49 == reqIndex | way0V_73; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3669 = 7'h4a == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1365 = 7'h4a == reqIndex | way0V_74; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3670 = 7'h4b == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1366 = 7'h4b == reqIndex | way0V_75; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3671 = 7'h4c == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1367 = 7'h4c == reqIndex | way0V_76; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3672 = 7'h4d == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1368 = 7'h4d == reqIndex | way0V_77; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3673 = 7'h4e == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1369 = 7'h4e == reqIndex | way0V_78; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3674 = 7'h4f == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1370 = 7'h4f == reqIndex | way0V_79; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3675 = 7'h50 == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1371 = 7'h50 == reqIndex | way0V_80; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3676 = 7'h51 == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1372 = 7'h51 == reqIndex | way0V_81; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3677 = 7'h52 == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1373 = 7'h52 == reqIndex | way0V_82; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3678 = 7'h53 == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1374 = 7'h53 == reqIndex | way0V_83; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3679 = 7'h54 == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1375 = 7'h54 == reqIndex | way0V_84; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3680 = 7'h55 == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1376 = 7'h55 == reqIndex | way0V_85; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3681 = 7'h56 == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1377 = 7'h56 == reqIndex | way0V_86; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3682 = 7'h57 == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1378 = 7'h57 == reqIndex | way0V_87; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3683 = 7'h58 == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1379 = 7'h58 == reqIndex | way0V_88; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3684 = 7'h59 == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1380 = 7'h59 == reqIndex | way0V_89; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3685 = 7'h5a == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1381 = 7'h5a == reqIndex | way0V_90; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3686 = 7'h5b == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1382 = 7'h5b == reqIndex | way0V_91; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3687 = 7'h5c == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1383 = 7'h5c == reqIndex | way0V_92; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3688 = 7'h5d == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1384 = 7'h5d == reqIndex | way0V_93; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3689 = 7'h5e == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1385 = 7'h5e == reqIndex | way0V_94; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3690 = 7'h5f == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1386 = 7'h5f == reqIndex | way0V_95; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3691 = 7'h60 == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1387 = 7'h60 == reqIndex | way0V_96; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3692 = 7'h61 == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1388 = 7'h61 == reqIndex | way0V_97; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3693 = 7'h62 == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1389 = 7'h62 == reqIndex | way0V_98; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3694 = 7'h63 == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1390 = 7'h63 == reqIndex | way0V_99; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3695 = 7'h64 == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1391 = 7'h64 == reqIndex | way0V_100; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3696 = 7'h65 == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1392 = 7'h65 == reqIndex | way0V_101; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3697 = 7'h66 == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1393 = 7'h66 == reqIndex | way0V_102; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3698 = 7'h67 == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1394 = 7'h67 == reqIndex | way0V_103; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3699 = 7'h68 == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1395 = 7'h68 == reqIndex | way0V_104; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3700 = 7'h69 == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1396 = 7'h69 == reqIndex | way0V_105; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3701 = 7'h6a == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1397 = 7'h6a == reqIndex | way0V_106; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3702 = 7'h6b == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1398 = 7'h6b == reqIndex | way0V_107; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3703 = 7'h6c == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1399 = 7'h6c == reqIndex | way0V_108; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3704 = 7'h6d == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1400 = 7'h6d == reqIndex | way0V_109; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3705 = 7'h6e == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1401 = 7'h6e == reqIndex | way0V_110; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3706 = 7'h6f == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1402 = 7'h6f == reqIndex | way0V_111; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3707 = 7'h70 == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1403 = 7'h70 == reqIndex | way0V_112; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3708 = 7'h71 == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1404 = 7'h71 == reqIndex | way0V_113; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3709 = 7'h72 == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1405 = 7'h72 == reqIndex | way0V_114; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3710 = 7'h73 == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1406 = 7'h73 == reqIndex | way0V_115; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3711 = 7'h74 == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1407 = 7'h74 == reqIndex | way0V_116; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3712 = 7'h75 == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1408 = 7'h75 == reqIndex | way0V_117; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3713 = 7'h76 == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1409 = 7'h76 == reqIndex | way0V_118; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3714 = 7'h77 == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1410 = 7'h77 == reqIndex | way0V_119; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3715 = 7'h78 == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1411 = 7'h78 == reqIndex | way0V_120; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3716 = 7'h79 == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1412 = 7'h79 == reqIndex | way0V_121; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3717 = 7'h7a == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1413 = 7'h7a == reqIndex | way0V_122; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3718 = 7'h7b == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1414 = 7'h7b == reqIndex | way0V_123; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3719 = 7'h7c == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1415 = 7'h7c == reqIndex | way0V_124; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3720 = 7'h7d == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1416 = 7'h7d == reqIndex | way0V_125; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3721 = 7'h7e == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1417 = 7'h7e == reqIndex | way0V_126; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_3722 = 7'h7f == reqIndex; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1418 = 7'h7f == reqIndex | way0V_127; // @[DCache.scala 177:{23,23} 33:22]
  wire  _GEN_1675 = _GEN_3595 | way1V_0; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1676 = _GEN_3596 | way1V_1; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1677 = _GEN_3597 | way1V_2; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1678 = _GEN_3598 | way1V_3; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1679 = _GEN_3599 | way1V_4; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1680 = _GEN_3600 | way1V_5; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1681 = _GEN_3601 | way1V_6; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1682 = _GEN_3602 | way1V_7; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1683 = _GEN_3603 | way1V_8; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1684 = _GEN_3604 | way1V_9; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1685 = _GEN_3605 | way1V_10; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1686 = _GEN_3606 | way1V_11; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1687 = _GEN_3607 | way1V_12; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1688 = _GEN_3608 | way1V_13; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1689 = _GEN_3609 | way1V_14; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1690 = _GEN_3610 | way1V_15; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1691 = _GEN_3611 | way1V_16; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1692 = _GEN_3612 | way1V_17; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1693 = _GEN_3613 | way1V_18; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1694 = _GEN_3614 | way1V_19; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1695 = _GEN_3615 | way1V_20; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1696 = _GEN_3616 | way1V_21; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1697 = _GEN_3617 | way1V_22; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1698 = _GEN_3618 | way1V_23; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1699 = _GEN_3619 | way1V_24; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1700 = _GEN_3620 | way1V_25; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1701 = _GEN_3621 | way1V_26; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1702 = _GEN_3622 | way1V_27; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1703 = _GEN_3623 | way1V_28; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1704 = _GEN_3624 | way1V_29; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1705 = _GEN_3625 | way1V_30; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1706 = _GEN_3626 | way1V_31; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1707 = _GEN_3627 | way1V_32; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1708 = _GEN_3628 | way1V_33; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1709 = _GEN_3629 | way1V_34; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1710 = _GEN_3630 | way1V_35; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1711 = _GEN_3631 | way1V_36; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1712 = _GEN_3632 | way1V_37; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1713 = _GEN_3633 | way1V_38; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1714 = _GEN_3634 | way1V_39; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1715 = _GEN_3635 | way1V_40; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1716 = _GEN_3636 | way1V_41; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1717 = _GEN_3637 | way1V_42; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1718 = _GEN_3638 | way1V_43; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1719 = _GEN_3639 | way1V_44; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1720 = _GEN_3640 | way1V_45; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1721 = _GEN_3641 | way1V_46; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1722 = _GEN_3642 | way1V_47; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1723 = _GEN_3643 | way1V_48; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1724 = _GEN_3644 | way1V_49; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1725 = _GEN_3645 | way1V_50; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1726 = _GEN_3646 | way1V_51; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1727 = _GEN_3647 | way1V_52; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1728 = _GEN_3648 | way1V_53; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1729 = _GEN_3649 | way1V_54; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1730 = _GEN_3650 | way1V_55; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1731 = _GEN_3651 | way1V_56; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1732 = _GEN_3652 | way1V_57; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1733 = _GEN_3653 | way1V_58; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1734 = _GEN_3654 | way1V_59; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1735 = _GEN_3655 | way1V_60; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1736 = _GEN_3656 | way1V_61; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1737 = _GEN_3657 | way1V_62; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1738 = _GEN_3658 | way1V_63; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1739 = _GEN_3659 | way1V_64; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1740 = _GEN_3660 | way1V_65; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1741 = _GEN_3661 | way1V_66; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1742 = _GEN_3662 | way1V_67; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1743 = _GEN_3663 | way1V_68; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1744 = _GEN_3664 | way1V_69; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1745 = _GEN_3665 | way1V_70; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1746 = _GEN_3666 | way1V_71; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1747 = _GEN_3667 | way1V_72; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1748 = _GEN_3668 | way1V_73; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1749 = _GEN_3669 | way1V_74; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1750 = _GEN_3670 | way1V_75; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1751 = _GEN_3671 | way1V_76; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1752 = _GEN_3672 | way1V_77; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1753 = _GEN_3673 | way1V_78; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1754 = _GEN_3674 | way1V_79; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1755 = _GEN_3675 | way1V_80; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1756 = _GEN_3676 | way1V_81; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1757 = _GEN_3677 | way1V_82; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1758 = _GEN_3678 | way1V_83; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1759 = _GEN_3679 | way1V_84; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1760 = _GEN_3680 | way1V_85; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1761 = _GEN_3681 | way1V_86; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1762 = _GEN_3682 | way1V_87; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1763 = _GEN_3683 | way1V_88; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1764 = _GEN_3684 | way1V_89; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1765 = _GEN_3685 | way1V_90; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1766 = _GEN_3686 | way1V_91; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1767 = _GEN_3687 | way1V_92; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1768 = _GEN_3688 | way1V_93; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1769 = _GEN_3689 | way1V_94; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1770 = _GEN_3690 | way1V_95; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1771 = _GEN_3691 | way1V_96; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1772 = _GEN_3692 | way1V_97; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1773 = _GEN_3693 | way1V_98; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1774 = _GEN_3694 | way1V_99; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1775 = _GEN_3695 | way1V_100; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1776 = _GEN_3696 | way1V_101; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1777 = _GEN_3697 | way1V_102; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1778 = _GEN_3698 | way1V_103; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1779 = _GEN_3699 | way1V_104; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1780 = _GEN_3700 | way1V_105; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1781 = _GEN_3701 | way1V_106; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1782 = _GEN_3702 | way1V_107; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1783 = _GEN_3703 | way1V_108; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1784 = _GEN_3704 | way1V_109; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1785 = _GEN_3705 | way1V_110; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1786 = _GEN_3706 | way1V_111; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1787 = _GEN_3707 | way1V_112; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1788 = _GEN_3708 | way1V_113; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1789 = _GEN_3709 | way1V_114; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1790 = _GEN_3710 | way1V_115; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1791 = _GEN_3711 | way1V_116; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1792 = _GEN_3712 | way1V_117; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1793 = _GEN_3713 | way1V_118; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1794 = _GEN_3714 | way1V_119; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1795 = _GEN_3715 | way1V_120; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1796 = _GEN_3716 | way1V_121; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1797 = _GEN_3717 | way1V_122; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1798 = _GEN_3718 | way1V_123; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1799 = _GEN_3719 | way1V_124; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1800 = _GEN_3720 | way1V_125; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1801 = _GEN_3721 | way1V_126; // @[DCache.scala 181:{23,23} 39:22]
  wire  _GEN_1802 = _GEN_3722 | way1V_127; // @[DCache.scala 181:{23,23} 39:22]
  wire [127:0] _rData_T = sDoneEn ? io_out_data_read : 128'h0; // @[DCache.scala 188:20]
  wire [127:0] rData = sHitEn ? cacheRData : _rData_T; // @[DCache.scala 187:18]
  wire [63:0] rDataHL = reqOff[3] ? rData[127:64] : rData[63:0]; // @[DCache.scala 189:20]
  wire [8:0] _io_dmem_data_read_T_2 = {1'h0,rDataHL[7:0]}; // @[Cat.scala 31:58]
  wire [8:0] _io_dmem_data_read_T_4 = {1'h0,rDataHL[15:8]}; // @[Cat.scala 31:58]
  wire [8:0] _io_dmem_data_read_T_6 = {1'h0,rDataHL[23:16]}; // @[Cat.scala 31:58]
  wire [8:0] _io_dmem_data_read_T_8 = {1'h0,rDataHL[31:24]}; // @[Cat.scala 31:58]
  wire [8:0] _io_dmem_data_read_T_10 = {1'h0,rDataHL[39:32]}; // @[Cat.scala 31:58]
  wire [8:0] _io_dmem_data_read_T_12 = {1'h0,rDataHL[47:40]}; // @[Cat.scala 31:58]
  wire [8:0] _io_dmem_data_read_T_14 = {1'h0,rDataHL[55:48]}; // @[Cat.scala 31:58]
  wire [8:0] _io_dmem_data_read_T_16 = {1'h0,rDataHL[63:56]}; // @[Cat.scala 31:58]
  wire [8:0] _io_dmem_data_read_T_18 = 3'h1 == reqOff[2:0] ? _io_dmem_data_read_T_4 : _io_dmem_data_read_T_2; // @[Mux.scala 81:58]
  wire [8:0] _io_dmem_data_read_T_20 = 3'h2 == reqOff[2:0] ? _io_dmem_data_read_T_6 : _io_dmem_data_read_T_18; // @[Mux.scala 81:58]
  wire [8:0] _io_dmem_data_read_T_22 = 3'h3 == reqOff[2:0] ? _io_dmem_data_read_T_8 : _io_dmem_data_read_T_20; // @[Mux.scala 81:58]
  wire [8:0] _io_dmem_data_read_T_24 = 3'h4 == reqOff[2:0] ? _io_dmem_data_read_T_10 : _io_dmem_data_read_T_22; // @[Mux.scala 81:58]
  wire [8:0] _io_dmem_data_read_T_26 = 3'h5 == reqOff[2:0] ? _io_dmem_data_read_T_12 : _io_dmem_data_read_T_24; // @[Mux.scala 81:58]
  wire [8:0] _io_dmem_data_read_T_28 = 3'h6 == reqOff[2:0] ? _io_dmem_data_read_T_14 : _io_dmem_data_read_T_26; // @[Mux.scala 81:58]
  wire [8:0] _io_dmem_data_read_T_30 = 3'h7 == reqOff[2:0] ? _io_dmem_data_read_T_16 : _io_dmem_data_read_T_28; // @[Mux.scala 81:58]
  wire [16:0] _io_dmem_data_read_T_33 = {1'h0,rDataHL[15:0]}; // @[Cat.scala 31:58]
  wire [16:0] _io_dmem_data_read_T_35 = {1'h0,rDataHL[31:16]}; // @[Cat.scala 31:58]
  wire [16:0] _io_dmem_data_read_T_37 = {1'h0,rDataHL[47:32]}; // @[Cat.scala 31:58]
  wire [16:0] _io_dmem_data_read_T_39 = {1'h0,rDataHL[63:48]}; // @[Cat.scala 31:58]
  wire [16:0] _io_dmem_data_read_T_41 = 2'h1 == reqOff[2:1] ? _io_dmem_data_read_T_35 : _io_dmem_data_read_T_33; // @[Mux.scala 81:58]
  wire [16:0] _io_dmem_data_read_T_43 = 2'h2 == reqOff[2:1] ? _io_dmem_data_read_T_37 : _io_dmem_data_read_T_41; // @[Mux.scala 81:58]
  wire [16:0] _io_dmem_data_read_T_45 = 2'h3 == reqOff[2:1] ? _io_dmem_data_read_T_39 : _io_dmem_data_read_T_43; // @[Mux.scala 81:58]
  wire [32:0] _io_dmem_data_read_T_48 = {1'h0,rDataHL[31:0]}; // @[Cat.scala 31:58]
  wire [32:0] _io_dmem_data_read_T_50 = {1'h0,rDataHL[63:32]}; // @[Cat.scala 31:58]
  wire [32:0] _io_dmem_data_read_T_52 = reqOff[2] ? _io_dmem_data_read_T_50 : _io_dmem_data_read_T_48; // @[Mux.scala 81:58]
  wire [16:0] _io_dmem_data_read_T_54 = 2'h1 == io_dmem_data_size ? _io_dmem_data_read_T_45 : {{8'd0},
    _io_dmem_data_read_T_30}; // @[Mux.scala 81:58]
  wire [32:0] _io_dmem_data_read_T_56 = 2'h2 == io_dmem_data_size ? _io_dmem_data_read_T_52 : {{16'd0},
    _io_dmem_data_read_T_54}; // @[Mux.scala 81:58]
  wire  cacheIndex = _cacheIndex_T_3[0];
  S011HD1P_X32Y2D128_BW req ( // @[DCache.scala 225:19]
    .Q(req_Q),
    .CLK(req_CLK),
    .CEN(req_CEN),
    .WEN(req_WEN),
    .BWEN(req_BWEN),
    .A(req_A),
    .D(req_D)
  );
  assign io_dmem_data_ready = sHitEn & cacheHitEn | sDoneEn; // @[DCache.scala 191:43]
  assign io_dmem_data_read = 2'h3 == io_dmem_data_size ? rDataHL : {{31'd0}, _io_dmem_data_read_T_56}; // @[Mux.scala 81:58]
  assign io_out_data_valid = sWriteEn | sCacheWEn; // @[DCache.scala 216:24]
  assign io_out_data_req = state == 3'h3; // @[DCache.scala 134:24]
  assign io_out_data_addr = io_dmem_data_addr; // @[DCache.scala 219:17]
  assign io_out_data_strb = sWriteEn ? io_dmem_data_strb : 8'h0; // @[DCache.scala 221:23]
  assign io_out_data_write = sWriteEn ? cacheRData : 128'h0; // @[DCache.scala 222:24]
  assign req_CLK = clock; // @[DCache.scala 226:14]
  assign req_CEN = 1'h1; // @[DCache.scala 227:14]
  assign req_WEN = io_dmem_data_req ? cacheHitEn : sCacheWEn; // @[DCache.scala 168:19]
  assign req_BWEN = io_dmem_data_req ? {{63'd0}, valid_strb} : 128'hffffffffffffffffffffffffffffffff; // @[DCache.scala 170:20]
  assign req_A = {{7'd0}, cacheIndex}; // @[DCache.scala 231:12]
  assign req_D = _valid_WData_T[127:0]; // @[DCache.scala 232:12]
  always @(posedge clock) begin
    if (reset) begin // @[DCache.scala 33:22]
      way0V_0 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_0 <= _GEN_1291;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_1 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_1 <= _GEN_1292;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_2 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_2 <= _GEN_1293;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_3 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_3 <= _GEN_1294;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_4 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_4 <= _GEN_1295;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_5 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_5 <= _GEN_1296;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_6 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_6 <= _GEN_1297;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_7 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_7 <= _GEN_1298;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_8 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_8 <= _GEN_1299;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_9 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_9 <= _GEN_1300;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_10 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_10 <= _GEN_1301;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_11 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_11 <= _GEN_1302;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_12 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_12 <= _GEN_1303;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_13 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_13 <= _GEN_1304;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_14 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_14 <= _GEN_1305;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_15 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_15 <= _GEN_1306;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_16 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_16 <= _GEN_1307;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_17 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_17 <= _GEN_1308;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_18 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_18 <= _GEN_1309;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_19 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_19 <= _GEN_1310;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_20 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_20 <= _GEN_1311;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_21 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_21 <= _GEN_1312;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_22 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_22 <= _GEN_1313;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_23 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_23 <= _GEN_1314;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_24 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_24 <= _GEN_1315;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_25 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_25 <= _GEN_1316;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_26 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_26 <= _GEN_1317;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_27 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_27 <= _GEN_1318;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_28 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_28 <= _GEN_1319;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_29 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_29 <= _GEN_1320;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_30 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_30 <= _GEN_1321;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_31 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_31 <= _GEN_1322;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_32 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_32 <= _GEN_1323;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_33 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_33 <= _GEN_1324;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_34 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_34 <= _GEN_1325;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_35 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_35 <= _GEN_1326;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_36 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_36 <= _GEN_1327;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_37 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_37 <= _GEN_1328;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_38 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_38 <= _GEN_1329;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_39 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_39 <= _GEN_1330;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_40 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_40 <= _GEN_1331;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_41 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_41 <= _GEN_1332;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_42 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_42 <= _GEN_1333;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_43 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_43 <= _GEN_1334;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_44 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_44 <= _GEN_1335;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_45 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_45 <= _GEN_1336;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_46 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_46 <= _GEN_1337;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_47 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_47 <= _GEN_1338;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_48 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_48 <= _GEN_1339;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_49 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_49 <= _GEN_1340;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_50 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_50 <= _GEN_1341;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_51 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_51 <= _GEN_1342;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_52 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_52 <= _GEN_1343;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_53 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_53 <= _GEN_1344;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_54 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_54 <= _GEN_1345;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_55 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_55 <= _GEN_1346;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_56 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_56 <= _GEN_1347;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_57 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_57 <= _GEN_1348;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_58 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_58 <= _GEN_1349;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_59 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_59 <= _GEN_1350;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_60 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_60 <= _GEN_1351;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_61 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_61 <= _GEN_1352;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_62 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_62 <= _GEN_1353;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_63 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_63 <= _GEN_1354;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_64 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_64 <= _GEN_1355;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_65 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_65 <= _GEN_1356;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_66 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_66 <= _GEN_1357;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_67 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_67 <= _GEN_1358;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_68 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_68 <= _GEN_1359;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_69 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_69 <= _GEN_1360;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_70 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_70 <= _GEN_1361;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_71 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_71 <= _GEN_1362;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_72 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_72 <= _GEN_1363;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_73 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_73 <= _GEN_1364;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_74 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_74 <= _GEN_1365;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_75 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_75 <= _GEN_1366;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_76 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_76 <= _GEN_1367;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_77 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_77 <= _GEN_1368;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_78 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_78 <= _GEN_1369;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_79 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_79 <= _GEN_1370;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_80 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_80 <= _GEN_1371;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_81 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_81 <= _GEN_1372;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_82 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_82 <= _GEN_1373;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_83 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_83 <= _GEN_1374;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_84 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_84 <= _GEN_1375;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_85 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_85 <= _GEN_1376;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_86 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_86 <= _GEN_1377;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_87 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_87 <= _GEN_1378;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_88 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_88 <= _GEN_1379;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_89 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_89 <= _GEN_1380;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_90 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_90 <= _GEN_1381;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_91 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_91 <= _GEN_1382;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_92 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_92 <= _GEN_1383;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_93 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_93 <= _GEN_1384;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_94 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_94 <= _GEN_1385;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_95 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_95 <= _GEN_1386;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_96 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_96 <= _GEN_1387;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_97 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_97 <= _GEN_1388;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_98 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_98 <= _GEN_1389;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_99 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_99 <= _GEN_1390;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_100 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_100 <= _GEN_1391;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_101 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_101 <= _GEN_1392;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_102 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_102 <= _GEN_1393;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_103 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_103 <= _GEN_1394;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_104 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_104 <= _GEN_1395;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_105 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_105 <= _GEN_1396;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_106 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_106 <= _GEN_1397;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_107 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_107 <= _GEN_1398;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_108 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_108 <= _GEN_1399;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_109 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_109 <= _GEN_1400;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_110 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_110 <= _GEN_1401;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_111 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_111 <= _GEN_1402;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_112 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_112 <= _GEN_1403;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_113 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_113 <= _GEN_1404;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_114 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_114 <= _GEN_1405;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_115 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_115 <= _GEN_1406;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_116 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_116 <= _GEN_1407;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_117 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_117 <= _GEN_1408;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_118 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_118 <= _GEN_1409;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_119 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_119 <= _GEN_1410;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_120 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_120 <= _GEN_1411;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_121 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_121 <= _GEN_1412;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_122 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_122 <= _GEN_1413;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_123 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_123 <= _GEN_1414;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_124 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_124 <= _GEN_1415;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_125 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_125 <= _GEN_1416;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_126 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_126 <= _GEN_1417;
      end
    end
    if (reset) begin // @[DCache.scala 33:22]
      way0V_127 <= 1'h0; // @[DCache.scala 33:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        way0V_127 <= _GEN_1418;
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_0 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h0 == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_0 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_1 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h1 == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_1 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_2 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h2 == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_2 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_3 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h3 == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_3 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_4 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h4 == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_4 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_5 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h5 == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_5 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_6 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h6 == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_6 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_7 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h7 == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_7 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_8 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h8 == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_8 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_9 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h9 == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_9 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_10 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'ha == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_10 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_11 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'hb == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_11 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_12 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'hc == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_12 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_13 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'hd == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_13 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_14 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'he == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_14 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_15 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'hf == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_15 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_16 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h10 == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_16 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_17 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h11 == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_17 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_18 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h12 == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_18 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_19 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h13 == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_19 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_20 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h14 == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_20 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_21 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h15 == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_21 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_22 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h16 == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_22 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_23 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h17 == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_23 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_24 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h18 == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_24 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_25 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h19 == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_25 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_26 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h1a == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_26 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_27 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h1b == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_27 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_28 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h1c == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_28 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_29 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h1d == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_29 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_30 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h1e == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_30 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_31 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h1f == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_31 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_32 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h20 == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_32 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_33 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h21 == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_33 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_34 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h22 == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_34 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_35 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h23 == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_35 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_36 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h24 == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_36 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_37 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h25 == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_37 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_38 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h26 == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_38 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_39 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h27 == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_39 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_40 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h28 == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_40 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_41 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h29 == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_41 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_42 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h2a == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_42 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_43 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h2b == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_43 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_44 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h2c == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_44 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_45 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h2d == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_45 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_46 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h2e == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_46 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_47 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h2f == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_47 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_48 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h30 == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_48 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_49 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h31 == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_49 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_50 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h32 == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_50 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_51 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h33 == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_51 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_52 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h34 == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_52 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_53 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h35 == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_53 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_54 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h36 == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_54 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_55 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h37 == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_55 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_56 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h38 == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_56 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_57 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h39 == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_57 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_58 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h3a == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_58 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_59 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h3b == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_59 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_60 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h3c == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_60 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_61 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h3d == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_61 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_62 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h3e == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_62 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_63 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h3f == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_63 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_64 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h40 == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_64 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_65 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h41 == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_65 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_66 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h42 == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_66 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_67 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h43 == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_67 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_68 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h44 == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_68 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_69 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h45 == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_69 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_70 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h46 == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_70 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_71 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h47 == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_71 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_72 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h48 == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_72 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_73 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h49 == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_73 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_74 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h4a == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_74 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_75 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h4b == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_75 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_76 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h4c == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_76 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_77 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h4d == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_77 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_78 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h4e == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_78 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_79 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h4f == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_79 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_80 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h50 == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_80 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_81 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h51 == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_81 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_82 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h52 == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_82 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_83 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h53 == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_83 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_84 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h54 == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_84 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_85 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h55 == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_85 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_86 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h56 == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_86 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_87 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h57 == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_87 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_88 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h58 == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_88 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_89 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h59 == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_89 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_90 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h5a == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_90 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_91 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h5b == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_91 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_92 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h5c == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_92 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_93 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h5d == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_93 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_94 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h5e == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_94 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_95 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h5f == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_95 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_96 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h60 == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_96 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_97 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h61 == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_97 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_98 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h62 == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_98 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_99 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h63 == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_99 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_100 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h64 == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_100 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_101 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h65 == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_101 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_102 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h66 == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_102 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_103 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h67 == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_103 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_104 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h68 == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_104 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_105 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h69 == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_105 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_106 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h6a == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_106 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_107 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h6b == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_107 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_108 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h6c == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_108 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_109 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h6d == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_109 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_110 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h6e == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_110 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_111 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h6f == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_111 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_112 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h70 == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_112 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_113 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h71 == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_113 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_114 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h72 == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_114 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_115 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h73 == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_115 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_116 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h74 == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_116 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_117 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h75 == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_117 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_118 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h76 == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_118 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_119 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h77 == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_119 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_120 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h78 == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_120 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_121 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h79 == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_121 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_122 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h7a == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_122 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_123 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h7b == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_123 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_124 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h7c == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_124 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_125 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h7d == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_125 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_126 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h7e == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_126 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 34:24]
      way0Tag_127 <= 21'h0; // @[DCache.scala 34:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h7f == reqIndex) begin // @[DCache.scala 178:25]
          way0Tag_127 <= reqTag; // @[DCache.scala 178:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_0 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h0 == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_0 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_1 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h1 == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_1 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_2 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h2 == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_2 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_3 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h3 == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_3 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_4 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h4 == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_4 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_5 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h5 == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_5 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_6 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h6 == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_6 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_7 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h7 == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_7 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_8 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h8 == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_8 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_9 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h9 == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_9 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_10 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'ha == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_10 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_11 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'hb == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_11 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_12 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'hc == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_12 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_13 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'hd == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_13 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_14 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'he == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_14 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_15 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'hf == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_15 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_16 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h10 == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_16 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_17 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h11 == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_17 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_18 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h12 == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_18 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_19 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h13 == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_19 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_20 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h14 == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_20 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_21 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h15 == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_21 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_22 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h16 == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_22 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_23 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h17 == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_23 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_24 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h18 == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_24 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_25 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h19 == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_25 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_26 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h1a == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_26 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_27 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h1b == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_27 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_28 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h1c == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_28 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_29 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h1d == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_29 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_30 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h1e == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_30 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_31 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h1f == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_31 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_32 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h20 == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_32 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_33 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h21 == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_33 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_34 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h22 == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_34 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_35 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h23 == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_35 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_36 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h24 == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_36 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_37 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h25 == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_37 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_38 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h26 == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_38 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_39 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h27 == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_39 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_40 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h28 == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_40 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_41 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h29 == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_41 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_42 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h2a == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_42 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_43 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h2b == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_43 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_44 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h2c == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_44 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_45 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h2d == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_45 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_46 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h2e == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_46 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_47 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h2f == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_47 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_48 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h30 == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_48 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_49 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h31 == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_49 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_50 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h32 == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_50 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_51 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h33 == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_51 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_52 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h34 == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_52 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_53 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h35 == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_53 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_54 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h36 == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_54 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_55 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h37 == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_55 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_56 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h38 == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_56 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_57 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h39 == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_57 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_58 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h3a == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_58 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_59 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h3b == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_59 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_60 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h3c == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_60 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_61 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h3d == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_61 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_62 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h3e == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_62 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_63 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h3f == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_63 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_64 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h40 == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_64 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_65 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h41 == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_65 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_66 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h42 == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_66 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_67 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h43 == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_67 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_68 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h44 == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_68 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_69 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h45 == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_69 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_70 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h46 == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_70 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_71 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h47 == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_71 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_72 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h48 == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_72 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_73 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h49 == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_73 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_74 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h4a == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_74 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_75 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h4b == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_75 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_76 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h4c == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_76 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_77 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h4d == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_77 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_78 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h4e == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_78 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_79 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h4f == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_79 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_80 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h50 == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_80 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_81 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h51 == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_81 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_82 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h52 == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_82 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_83 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h53 == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_83 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_84 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h54 == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_84 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_85 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h55 == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_85 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_86 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h56 == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_86 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_87 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h57 == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_87 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_88 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h58 == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_88 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_89 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h59 == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_89 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_90 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h5a == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_90 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_91 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h5b == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_91 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_92 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h5c == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_92 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_93 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h5d == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_93 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_94 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h5e == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_94 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_95 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h5f == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_95 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_96 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h60 == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_96 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_97 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h61 == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_97 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_98 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h62 == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_98 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_99 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h63 == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_99 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_100 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h64 == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_100 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_101 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h65 == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_101 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_102 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h66 == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_102 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_103 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h67 == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_103 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_104 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h68 == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_104 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_105 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h69 == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_105 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_106 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h6a == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_106 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_107 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h6b == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_107 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_108 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h6c == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_108 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_109 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h6d == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_109 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_110 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h6e == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_110 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_111 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h6f == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_111 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_112 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h70 == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_112 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_113 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h71 == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_113 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_114 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h72 == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_114 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_115 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h73 == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_115 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_116 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h74 == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_116 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_117 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h75 == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_117 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_118 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h76 == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_118 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_119 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h77 == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_119 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_120 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h78 == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_120 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_121 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h79 == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_121 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_122 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h7a == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_122 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_123 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h7b == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_123 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_124 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h7c == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_124 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_125 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h7d == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_125 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_126 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h7e == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_126 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 36:24]
      way0Age_127 <= 1'h0; // @[DCache.scala 36:24]
    end else if (7'h7f == reqIndex) begin // @[DCache.scala 173:21]
      way0Age_127 <= ageWay0En & sDoneEn; // @[DCache.scala 173:21]
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_0 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h0 == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_0 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_1 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h1 == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_1 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_2 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h2 == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_2 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_3 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h3 == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_3 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_4 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h4 == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_4 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_5 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h5 == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_5 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_6 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h6 == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_6 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_7 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h7 == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_7 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_8 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h8 == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_8 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_9 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h9 == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_9 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_10 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'ha == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_10 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_11 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'hb == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_11 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_12 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'hc == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_12 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_13 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'hd == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_13 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_14 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'he == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_14 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_15 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'hf == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_15 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_16 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h10 == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_16 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_17 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h11 == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_17 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_18 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h12 == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_18 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_19 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h13 == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_19 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_20 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h14 == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_20 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_21 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h15 == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_21 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_22 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h16 == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_22 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_23 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h17 == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_23 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_24 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h18 == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_24 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_25 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h19 == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_25 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_26 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h1a == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_26 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_27 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h1b == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_27 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_28 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h1c == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_28 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_29 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h1d == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_29 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_30 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h1e == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_30 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_31 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h1f == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_31 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_32 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h20 == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_32 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_33 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h21 == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_33 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_34 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h22 == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_34 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_35 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h23 == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_35 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_36 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h24 == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_36 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_37 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h25 == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_37 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_38 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h26 == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_38 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_39 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h27 == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_39 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_40 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h28 == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_40 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_41 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h29 == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_41 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_42 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h2a == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_42 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_43 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h2b == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_43 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_44 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h2c == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_44 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_45 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h2d == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_45 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_46 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h2e == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_46 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_47 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h2f == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_47 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_48 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h30 == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_48 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_49 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h31 == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_49 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_50 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h32 == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_50 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_51 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h33 == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_51 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_52 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h34 == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_52 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_53 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h35 == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_53 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_54 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h36 == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_54 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_55 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h37 == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_55 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_56 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h38 == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_56 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_57 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h39 == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_57 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_58 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h3a == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_58 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_59 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h3b == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_59 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_60 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h3c == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_60 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_61 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h3d == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_61 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_62 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h3e == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_62 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_63 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h3f == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_63 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_64 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h40 == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_64 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_65 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h41 == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_65 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_66 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h42 == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_66 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_67 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h43 == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_67 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_68 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h44 == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_68 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_69 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h45 == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_69 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_70 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h46 == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_70 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_71 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h47 == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_71 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_72 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h48 == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_72 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_73 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h49 == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_73 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_74 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h4a == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_74 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_75 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h4b == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_75 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_76 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h4c == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_76 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_77 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h4d == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_77 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_78 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h4e == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_78 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_79 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h4f == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_79 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_80 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h50 == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_80 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_81 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h51 == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_81 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_82 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h52 == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_82 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_83 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h53 == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_83 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_84 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h54 == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_84 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_85 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h55 == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_85 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_86 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h56 == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_86 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_87 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h57 == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_87 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_88 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h58 == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_88 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_89 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h59 == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_89 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_90 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h5a == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_90 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_91 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h5b == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_91 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_92 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h5c == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_92 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_93 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h5d == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_93 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_94 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h5e == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_94 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_95 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h5f == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_95 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_96 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h60 == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_96 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_97 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h61 == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_97 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_98 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h62 == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_98 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_99 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h63 == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_99 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_100 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h64 == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_100 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_101 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h65 == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_101 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_102 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h66 == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_102 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_103 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h67 == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_103 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_104 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h68 == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_104 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_105 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h69 == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_105 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_106 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h6a == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_106 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_107 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h6b == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_107 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_108 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h6c == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_108 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_109 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h6d == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_109 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_110 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h6e == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_110 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_111 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h6f == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_111 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_112 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h70 == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_112 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_113 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h71 == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_113 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_114 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h72 == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_114 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_115 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h73 == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_115 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_116 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h74 == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_116 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_117 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h75 == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_117 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_118 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h76 == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_118 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_119 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h77 == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_119 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_120 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h78 == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_120 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_121 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h79 == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_121 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_122 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h7a == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_122 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_123 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h7b == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_123 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_124 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h7c == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_124 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_125 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h7d == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_125 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_126 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h7e == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_126 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_127 <= 1'h0; // @[DCache.scala 37:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (cacheLineWay) begin // @[DCache.scala 176:24]
        if (7'h7f == reqIndex) begin // @[DCache.scala 179:27]
          way0Dirty_127 <= io_dmem_data_req; // @[DCache.scala 179:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_0 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_0 <= _GEN_1675;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_1 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_1 <= _GEN_1676;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_2 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_2 <= _GEN_1677;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_3 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_3 <= _GEN_1678;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_4 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_4 <= _GEN_1679;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_5 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_5 <= _GEN_1680;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_6 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_6 <= _GEN_1681;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_7 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_7 <= _GEN_1682;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_8 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_8 <= _GEN_1683;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_9 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_9 <= _GEN_1684;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_10 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_10 <= _GEN_1685;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_11 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_11 <= _GEN_1686;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_12 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_12 <= _GEN_1687;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_13 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_13 <= _GEN_1688;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_14 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_14 <= _GEN_1689;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_15 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_15 <= _GEN_1690;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_16 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_16 <= _GEN_1691;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_17 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_17 <= _GEN_1692;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_18 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_18 <= _GEN_1693;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_19 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_19 <= _GEN_1694;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_20 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_20 <= _GEN_1695;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_21 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_21 <= _GEN_1696;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_22 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_22 <= _GEN_1697;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_23 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_23 <= _GEN_1698;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_24 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_24 <= _GEN_1699;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_25 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_25 <= _GEN_1700;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_26 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_26 <= _GEN_1701;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_27 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_27 <= _GEN_1702;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_28 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_28 <= _GEN_1703;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_29 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_29 <= _GEN_1704;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_30 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_30 <= _GEN_1705;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_31 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_31 <= _GEN_1706;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_32 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_32 <= _GEN_1707;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_33 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_33 <= _GEN_1708;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_34 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_34 <= _GEN_1709;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_35 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_35 <= _GEN_1710;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_36 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_36 <= _GEN_1711;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_37 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_37 <= _GEN_1712;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_38 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_38 <= _GEN_1713;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_39 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_39 <= _GEN_1714;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_40 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_40 <= _GEN_1715;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_41 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_41 <= _GEN_1716;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_42 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_42 <= _GEN_1717;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_43 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_43 <= _GEN_1718;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_44 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_44 <= _GEN_1719;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_45 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_45 <= _GEN_1720;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_46 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_46 <= _GEN_1721;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_47 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_47 <= _GEN_1722;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_48 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_48 <= _GEN_1723;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_49 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_49 <= _GEN_1724;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_50 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_50 <= _GEN_1725;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_51 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_51 <= _GEN_1726;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_52 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_52 <= _GEN_1727;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_53 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_53 <= _GEN_1728;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_54 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_54 <= _GEN_1729;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_55 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_55 <= _GEN_1730;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_56 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_56 <= _GEN_1731;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_57 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_57 <= _GEN_1732;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_58 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_58 <= _GEN_1733;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_59 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_59 <= _GEN_1734;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_60 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_60 <= _GEN_1735;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_61 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_61 <= _GEN_1736;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_62 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_62 <= _GEN_1737;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_63 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_63 <= _GEN_1738;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_64 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_64 <= _GEN_1739;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_65 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_65 <= _GEN_1740;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_66 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_66 <= _GEN_1741;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_67 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_67 <= _GEN_1742;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_68 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_68 <= _GEN_1743;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_69 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_69 <= _GEN_1744;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_70 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_70 <= _GEN_1745;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_71 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_71 <= _GEN_1746;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_72 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_72 <= _GEN_1747;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_73 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_73 <= _GEN_1748;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_74 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_74 <= _GEN_1749;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_75 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_75 <= _GEN_1750;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_76 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_76 <= _GEN_1751;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_77 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_77 <= _GEN_1752;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_78 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_78 <= _GEN_1753;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_79 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_79 <= _GEN_1754;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_80 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_80 <= _GEN_1755;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_81 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_81 <= _GEN_1756;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_82 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_82 <= _GEN_1757;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_83 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_83 <= _GEN_1758;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_84 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_84 <= _GEN_1759;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_85 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_85 <= _GEN_1760;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_86 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_86 <= _GEN_1761;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_87 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_87 <= _GEN_1762;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_88 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_88 <= _GEN_1763;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_89 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_89 <= _GEN_1764;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_90 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_90 <= _GEN_1765;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_91 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_91 <= _GEN_1766;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_92 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_92 <= _GEN_1767;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_93 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_93 <= _GEN_1768;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_94 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_94 <= _GEN_1769;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_95 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_95 <= _GEN_1770;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_96 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_96 <= _GEN_1771;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_97 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_97 <= _GEN_1772;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_98 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_98 <= _GEN_1773;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_99 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_99 <= _GEN_1774;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_100 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_100 <= _GEN_1775;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_101 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_101 <= _GEN_1776;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_102 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_102 <= _GEN_1777;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_103 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_103 <= _GEN_1778;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_104 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_104 <= _GEN_1779;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_105 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_105 <= _GEN_1780;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_106 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_106 <= _GEN_1781;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_107 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_107 <= _GEN_1782;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_108 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_108 <= _GEN_1783;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_109 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_109 <= _GEN_1784;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_110 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_110 <= _GEN_1785;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_111 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_111 <= _GEN_1786;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_112 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_112 <= _GEN_1787;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_113 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_113 <= _GEN_1788;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_114 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_114 <= _GEN_1789;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_115 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_115 <= _GEN_1790;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_116 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_116 <= _GEN_1791;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_117 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_117 <= _GEN_1792;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_118 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_118 <= _GEN_1793;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_119 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_119 <= _GEN_1794;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_120 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_120 <= _GEN_1795;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_121 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_121 <= _GEN_1796;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_122 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_122 <= _GEN_1797;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_123 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_123 <= _GEN_1798;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_124 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_124 <= _GEN_1799;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_125 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_125 <= _GEN_1800;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_126 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_126 <= _GEN_1801;
      end
    end
    if (reset) begin // @[DCache.scala 39:22]
      way1V_127 <= 1'h0; // @[DCache.scala 39:22]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        way1V_127 <= _GEN_1802;
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_0 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h0 == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_0 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_1 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h1 == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_1 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_2 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h2 == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_2 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_3 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h3 == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_3 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_4 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h4 == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_4 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_5 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h5 == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_5 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_6 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h6 == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_6 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_7 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h7 == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_7 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_8 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h8 == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_8 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_9 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h9 == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_9 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_10 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'ha == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_10 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_11 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'hb == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_11 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_12 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'hc == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_12 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_13 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'hd == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_13 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_14 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'he == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_14 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_15 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'hf == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_15 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_16 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h10 == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_16 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_17 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h11 == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_17 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_18 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h12 == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_18 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_19 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h13 == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_19 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_20 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h14 == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_20 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_21 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h15 == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_21 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_22 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h16 == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_22 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_23 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h17 == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_23 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_24 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h18 == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_24 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_25 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h19 == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_25 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_26 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h1a == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_26 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_27 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h1b == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_27 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_28 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h1c == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_28 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_29 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h1d == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_29 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_30 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h1e == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_30 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_31 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h1f == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_31 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_32 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h20 == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_32 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_33 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h21 == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_33 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_34 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h22 == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_34 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_35 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h23 == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_35 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_36 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h24 == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_36 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_37 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h25 == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_37 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_38 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h26 == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_38 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_39 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h27 == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_39 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_40 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h28 == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_40 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_41 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h29 == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_41 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_42 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h2a == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_42 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_43 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h2b == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_43 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_44 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h2c == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_44 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_45 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h2d == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_45 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_46 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h2e == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_46 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_47 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h2f == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_47 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_48 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h30 == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_48 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_49 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h31 == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_49 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_50 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h32 == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_50 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_51 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h33 == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_51 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_52 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h34 == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_52 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_53 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h35 == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_53 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_54 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h36 == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_54 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_55 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h37 == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_55 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_56 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h38 == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_56 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_57 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h39 == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_57 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_58 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h3a == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_58 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_59 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h3b == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_59 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_60 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h3c == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_60 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_61 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h3d == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_61 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_62 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h3e == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_62 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_63 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h3f == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_63 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_64 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h40 == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_64 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_65 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h41 == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_65 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_66 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h42 == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_66 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_67 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h43 == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_67 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_68 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h44 == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_68 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_69 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h45 == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_69 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_70 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h46 == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_70 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_71 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h47 == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_71 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_72 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h48 == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_72 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_73 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h49 == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_73 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_74 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h4a == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_74 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_75 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h4b == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_75 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_76 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h4c == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_76 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_77 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h4d == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_77 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_78 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h4e == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_78 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_79 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h4f == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_79 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_80 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h50 == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_80 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_81 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h51 == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_81 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_82 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h52 == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_82 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_83 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h53 == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_83 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_84 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h54 == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_84 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_85 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h55 == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_85 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_86 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h56 == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_86 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_87 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h57 == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_87 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_88 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h58 == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_88 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_89 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h59 == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_89 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_90 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h5a == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_90 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_91 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h5b == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_91 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_92 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h5c == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_92 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_93 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h5d == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_93 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_94 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h5e == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_94 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_95 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h5f == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_95 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_96 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h60 == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_96 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_97 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h61 == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_97 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_98 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h62 == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_98 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_99 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h63 == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_99 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_100 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h64 == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_100 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_101 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h65 == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_101 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_102 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h66 == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_102 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_103 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h67 == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_103 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_104 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h68 == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_104 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_105 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h69 == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_105 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_106 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h6a == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_106 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_107 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h6b == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_107 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_108 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h6c == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_108 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_109 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h6d == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_109 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_110 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h6e == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_110 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_111 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h6f == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_111 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_112 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h70 == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_112 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_113 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h71 == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_113 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_114 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h72 == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_114 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_115 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h73 == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_115 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_116 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h74 == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_116 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_117 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h75 == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_117 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_118 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h76 == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_118 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_119 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h77 == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_119 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_120 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h78 == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_120 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_121 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h79 == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_121 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_122 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h7a == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_122 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_123 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h7b == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_123 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_124 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h7c == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_124 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_125 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h7d == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_125 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_126 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h7e == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_126 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:24]
      way1Tag_127 <= 21'h0; // @[DCache.scala 40:24]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h7f == reqIndex) begin // @[DCache.scala 182:25]
          way1Tag_127 <= reqTag; // @[DCache.scala 182:25]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_0 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h0 == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_0 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_1 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h1 == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_1 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_2 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h2 == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_2 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_3 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h3 == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_3 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_4 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h4 == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_4 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_5 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h5 == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_5 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_6 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h6 == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_6 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_7 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h7 == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_7 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_8 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h8 == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_8 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_9 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h9 == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_9 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_10 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'ha == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_10 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_11 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'hb == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_11 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_12 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'hc == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_12 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_13 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'hd == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_13 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_14 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'he == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_14 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_15 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'hf == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_15 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_16 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h10 == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_16 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_17 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h11 == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_17 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_18 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h12 == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_18 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_19 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h13 == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_19 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_20 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h14 == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_20 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_21 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h15 == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_21 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_22 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h16 == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_22 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_23 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h17 == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_23 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_24 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h18 == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_24 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_25 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h19 == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_25 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_26 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h1a == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_26 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_27 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h1b == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_27 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_28 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h1c == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_28 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_29 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h1d == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_29 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_30 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h1e == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_30 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_31 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h1f == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_31 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_32 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h20 == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_32 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_33 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h21 == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_33 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_34 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h22 == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_34 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_35 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h23 == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_35 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_36 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h24 == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_36 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_37 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h25 == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_37 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_38 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h26 == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_38 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_39 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h27 == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_39 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_40 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h28 == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_40 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_41 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h29 == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_41 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_42 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h2a == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_42 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_43 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h2b == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_43 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_44 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h2c == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_44 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_45 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h2d == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_45 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_46 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h2e == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_46 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_47 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h2f == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_47 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_48 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h30 == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_48 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_49 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h31 == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_49 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_50 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h32 == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_50 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_51 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h33 == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_51 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_52 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h34 == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_52 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_53 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h35 == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_53 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_54 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h36 == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_54 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_55 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h37 == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_55 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_56 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h38 == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_56 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_57 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h39 == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_57 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_58 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h3a == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_58 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_59 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h3b == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_59 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_60 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h3c == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_60 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_61 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h3d == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_61 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_62 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h3e == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_62 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_63 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h3f == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_63 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_64 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h40 == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_64 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_65 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h41 == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_65 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_66 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h42 == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_66 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_67 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h43 == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_67 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_68 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h44 == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_68 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_69 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h45 == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_69 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_70 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h46 == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_70 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_71 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h47 == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_71 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_72 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h48 == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_72 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_73 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h49 == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_73 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_74 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h4a == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_74 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_75 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h4b == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_75 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_76 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h4c == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_76 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_77 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h4d == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_77 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_78 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h4e == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_78 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_79 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h4f == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_79 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_80 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h50 == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_80 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_81 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h51 == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_81 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_82 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h52 == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_82 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_83 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h53 == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_83 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_84 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h54 == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_84 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_85 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h55 == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_85 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_86 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h56 == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_86 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_87 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h57 == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_87 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_88 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h58 == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_88 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_89 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h59 == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_89 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_90 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h5a == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_90 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_91 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h5b == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_91 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_92 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h5c == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_92 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_93 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h5d == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_93 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_94 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h5e == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_94 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_95 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h5f == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_95 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_96 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h60 == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_96 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_97 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h61 == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_97 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_98 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h62 == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_98 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_99 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h63 == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_99 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_100 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h64 == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_100 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_101 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h65 == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_101 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_102 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h66 == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_102 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_103 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h67 == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_103 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_104 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h68 == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_104 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_105 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h69 == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_105 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_106 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h6a == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_106 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_107 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h6b == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_107 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_108 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h6c == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_108 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_109 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h6d == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_109 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_110 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h6e == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_110 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_111 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h6f == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_111 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_112 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h70 == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_112 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_113 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h71 == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_113 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_114 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h72 == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_114 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_115 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h73 == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_115 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_116 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h74 == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_116 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_117 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h75 == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_117 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_118 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h76 == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_118 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_119 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h77 == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_119 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_120 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h78 == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_120 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_121 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h79 == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_121 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_122 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h7a == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_122 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_123 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h7b == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_123 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_124 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h7c == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_124 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_125 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h7d == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_125 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_126 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h7e == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_126 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_127 <= 1'h0; // @[DCache.scala 43:26]
    end else if (sDoneEn) begin // @[DCache.scala 175:17]
      if (!(cacheLineWay)) begin // @[DCache.scala 176:24]
        if (7'h7f == reqIndex) begin // @[DCache.scala 183:27]
          way1Dirty_127 <= io_dmem_data_req; // @[DCache.scala 183:27]
        end
      end
    end
    if (reset) begin // @[DCache.scala 46:22]
      state <= 3'h0; // @[DCache.scala 46:22]
    end else if (3'h0 == state) begin // @[DCache.scala 81:17]
      if (io_dmem_data_valid) begin // @[DCache.scala 83:29]
        state <= 3'h1; // @[DCache.scala 84:15]
      end
    end else if (3'h1 == state) begin // @[DCache.scala 81:17]
      if (cacheHitEn) begin // @[DCache.scala 88:27]
        state <= 3'h0; // @[DCache.scala 89:15]
      end else begin
        state <= 3'h2; // @[DCache.scala 91:15]
      end
    end else if (3'h2 == state) begin // @[DCache.scala 81:17]
      state <= _GEN_2;
    end else begin
      state <= _GEN_7;
    end
    cacheWriteEn_REG <= io_out_data_ready; // @[DCache.scala 164:41]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  way0V_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  way0V_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  way0V_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  way0V_3 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  way0V_4 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  way0V_5 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  way0V_6 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  way0V_7 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  way0V_8 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  way0V_9 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  way0V_10 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  way0V_11 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  way0V_12 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  way0V_13 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  way0V_14 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  way0V_15 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  way0V_16 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  way0V_17 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  way0V_18 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  way0V_19 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  way0V_20 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  way0V_21 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  way0V_22 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  way0V_23 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  way0V_24 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  way0V_25 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  way0V_26 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  way0V_27 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  way0V_28 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  way0V_29 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  way0V_30 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  way0V_31 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  way0V_32 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  way0V_33 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  way0V_34 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  way0V_35 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  way0V_36 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  way0V_37 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  way0V_38 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  way0V_39 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  way0V_40 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  way0V_41 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  way0V_42 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  way0V_43 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  way0V_44 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  way0V_45 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  way0V_46 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  way0V_47 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  way0V_48 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  way0V_49 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  way0V_50 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  way0V_51 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  way0V_52 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  way0V_53 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  way0V_54 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  way0V_55 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  way0V_56 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  way0V_57 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  way0V_58 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  way0V_59 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  way0V_60 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  way0V_61 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  way0V_62 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  way0V_63 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  way0V_64 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  way0V_65 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  way0V_66 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  way0V_67 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  way0V_68 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  way0V_69 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  way0V_70 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  way0V_71 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  way0V_72 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  way0V_73 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  way0V_74 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  way0V_75 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  way0V_76 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  way0V_77 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  way0V_78 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  way0V_79 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  way0V_80 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  way0V_81 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  way0V_82 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  way0V_83 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  way0V_84 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  way0V_85 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  way0V_86 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  way0V_87 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  way0V_88 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  way0V_89 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  way0V_90 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  way0V_91 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  way0V_92 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  way0V_93 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  way0V_94 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  way0V_95 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  way0V_96 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  way0V_97 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  way0V_98 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  way0V_99 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  way0V_100 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  way0V_101 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  way0V_102 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  way0V_103 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  way0V_104 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  way0V_105 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  way0V_106 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  way0V_107 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  way0V_108 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  way0V_109 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  way0V_110 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  way0V_111 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  way0V_112 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  way0V_113 = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  way0V_114 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  way0V_115 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  way0V_116 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  way0V_117 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  way0V_118 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  way0V_119 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  way0V_120 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  way0V_121 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  way0V_122 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  way0V_123 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  way0V_124 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  way0V_125 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  way0V_126 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  way0V_127 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  way0Tag_0 = _RAND_128[20:0];
  _RAND_129 = {1{`RANDOM}};
  way0Tag_1 = _RAND_129[20:0];
  _RAND_130 = {1{`RANDOM}};
  way0Tag_2 = _RAND_130[20:0];
  _RAND_131 = {1{`RANDOM}};
  way0Tag_3 = _RAND_131[20:0];
  _RAND_132 = {1{`RANDOM}};
  way0Tag_4 = _RAND_132[20:0];
  _RAND_133 = {1{`RANDOM}};
  way0Tag_5 = _RAND_133[20:0];
  _RAND_134 = {1{`RANDOM}};
  way0Tag_6 = _RAND_134[20:0];
  _RAND_135 = {1{`RANDOM}};
  way0Tag_7 = _RAND_135[20:0];
  _RAND_136 = {1{`RANDOM}};
  way0Tag_8 = _RAND_136[20:0];
  _RAND_137 = {1{`RANDOM}};
  way0Tag_9 = _RAND_137[20:0];
  _RAND_138 = {1{`RANDOM}};
  way0Tag_10 = _RAND_138[20:0];
  _RAND_139 = {1{`RANDOM}};
  way0Tag_11 = _RAND_139[20:0];
  _RAND_140 = {1{`RANDOM}};
  way0Tag_12 = _RAND_140[20:0];
  _RAND_141 = {1{`RANDOM}};
  way0Tag_13 = _RAND_141[20:0];
  _RAND_142 = {1{`RANDOM}};
  way0Tag_14 = _RAND_142[20:0];
  _RAND_143 = {1{`RANDOM}};
  way0Tag_15 = _RAND_143[20:0];
  _RAND_144 = {1{`RANDOM}};
  way0Tag_16 = _RAND_144[20:0];
  _RAND_145 = {1{`RANDOM}};
  way0Tag_17 = _RAND_145[20:0];
  _RAND_146 = {1{`RANDOM}};
  way0Tag_18 = _RAND_146[20:0];
  _RAND_147 = {1{`RANDOM}};
  way0Tag_19 = _RAND_147[20:0];
  _RAND_148 = {1{`RANDOM}};
  way0Tag_20 = _RAND_148[20:0];
  _RAND_149 = {1{`RANDOM}};
  way0Tag_21 = _RAND_149[20:0];
  _RAND_150 = {1{`RANDOM}};
  way0Tag_22 = _RAND_150[20:0];
  _RAND_151 = {1{`RANDOM}};
  way0Tag_23 = _RAND_151[20:0];
  _RAND_152 = {1{`RANDOM}};
  way0Tag_24 = _RAND_152[20:0];
  _RAND_153 = {1{`RANDOM}};
  way0Tag_25 = _RAND_153[20:0];
  _RAND_154 = {1{`RANDOM}};
  way0Tag_26 = _RAND_154[20:0];
  _RAND_155 = {1{`RANDOM}};
  way0Tag_27 = _RAND_155[20:0];
  _RAND_156 = {1{`RANDOM}};
  way0Tag_28 = _RAND_156[20:0];
  _RAND_157 = {1{`RANDOM}};
  way0Tag_29 = _RAND_157[20:0];
  _RAND_158 = {1{`RANDOM}};
  way0Tag_30 = _RAND_158[20:0];
  _RAND_159 = {1{`RANDOM}};
  way0Tag_31 = _RAND_159[20:0];
  _RAND_160 = {1{`RANDOM}};
  way0Tag_32 = _RAND_160[20:0];
  _RAND_161 = {1{`RANDOM}};
  way0Tag_33 = _RAND_161[20:0];
  _RAND_162 = {1{`RANDOM}};
  way0Tag_34 = _RAND_162[20:0];
  _RAND_163 = {1{`RANDOM}};
  way0Tag_35 = _RAND_163[20:0];
  _RAND_164 = {1{`RANDOM}};
  way0Tag_36 = _RAND_164[20:0];
  _RAND_165 = {1{`RANDOM}};
  way0Tag_37 = _RAND_165[20:0];
  _RAND_166 = {1{`RANDOM}};
  way0Tag_38 = _RAND_166[20:0];
  _RAND_167 = {1{`RANDOM}};
  way0Tag_39 = _RAND_167[20:0];
  _RAND_168 = {1{`RANDOM}};
  way0Tag_40 = _RAND_168[20:0];
  _RAND_169 = {1{`RANDOM}};
  way0Tag_41 = _RAND_169[20:0];
  _RAND_170 = {1{`RANDOM}};
  way0Tag_42 = _RAND_170[20:0];
  _RAND_171 = {1{`RANDOM}};
  way0Tag_43 = _RAND_171[20:0];
  _RAND_172 = {1{`RANDOM}};
  way0Tag_44 = _RAND_172[20:0];
  _RAND_173 = {1{`RANDOM}};
  way0Tag_45 = _RAND_173[20:0];
  _RAND_174 = {1{`RANDOM}};
  way0Tag_46 = _RAND_174[20:0];
  _RAND_175 = {1{`RANDOM}};
  way0Tag_47 = _RAND_175[20:0];
  _RAND_176 = {1{`RANDOM}};
  way0Tag_48 = _RAND_176[20:0];
  _RAND_177 = {1{`RANDOM}};
  way0Tag_49 = _RAND_177[20:0];
  _RAND_178 = {1{`RANDOM}};
  way0Tag_50 = _RAND_178[20:0];
  _RAND_179 = {1{`RANDOM}};
  way0Tag_51 = _RAND_179[20:0];
  _RAND_180 = {1{`RANDOM}};
  way0Tag_52 = _RAND_180[20:0];
  _RAND_181 = {1{`RANDOM}};
  way0Tag_53 = _RAND_181[20:0];
  _RAND_182 = {1{`RANDOM}};
  way0Tag_54 = _RAND_182[20:0];
  _RAND_183 = {1{`RANDOM}};
  way0Tag_55 = _RAND_183[20:0];
  _RAND_184 = {1{`RANDOM}};
  way0Tag_56 = _RAND_184[20:0];
  _RAND_185 = {1{`RANDOM}};
  way0Tag_57 = _RAND_185[20:0];
  _RAND_186 = {1{`RANDOM}};
  way0Tag_58 = _RAND_186[20:0];
  _RAND_187 = {1{`RANDOM}};
  way0Tag_59 = _RAND_187[20:0];
  _RAND_188 = {1{`RANDOM}};
  way0Tag_60 = _RAND_188[20:0];
  _RAND_189 = {1{`RANDOM}};
  way0Tag_61 = _RAND_189[20:0];
  _RAND_190 = {1{`RANDOM}};
  way0Tag_62 = _RAND_190[20:0];
  _RAND_191 = {1{`RANDOM}};
  way0Tag_63 = _RAND_191[20:0];
  _RAND_192 = {1{`RANDOM}};
  way0Tag_64 = _RAND_192[20:0];
  _RAND_193 = {1{`RANDOM}};
  way0Tag_65 = _RAND_193[20:0];
  _RAND_194 = {1{`RANDOM}};
  way0Tag_66 = _RAND_194[20:0];
  _RAND_195 = {1{`RANDOM}};
  way0Tag_67 = _RAND_195[20:0];
  _RAND_196 = {1{`RANDOM}};
  way0Tag_68 = _RAND_196[20:0];
  _RAND_197 = {1{`RANDOM}};
  way0Tag_69 = _RAND_197[20:0];
  _RAND_198 = {1{`RANDOM}};
  way0Tag_70 = _RAND_198[20:0];
  _RAND_199 = {1{`RANDOM}};
  way0Tag_71 = _RAND_199[20:0];
  _RAND_200 = {1{`RANDOM}};
  way0Tag_72 = _RAND_200[20:0];
  _RAND_201 = {1{`RANDOM}};
  way0Tag_73 = _RAND_201[20:0];
  _RAND_202 = {1{`RANDOM}};
  way0Tag_74 = _RAND_202[20:0];
  _RAND_203 = {1{`RANDOM}};
  way0Tag_75 = _RAND_203[20:0];
  _RAND_204 = {1{`RANDOM}};
  way0Tag_76 = _RAND_204[20:0];
  _RAND_205 = {1{`RANDOM}};
  way0Tag_77 = _RAND_205[20:0];
  _RAND_206 = {1{`RANDOM}};
  way0Tag_78 = _RAND_206[20:0];
  _RAND_207 = {1{`RANDOM}};
  way0Tag_79 = _RAND_207[20:0];
  _RAND_208 = {1{`RANDOM}};
  way0Tag_80 = _RAND_208[20:0];
  _RAND_209 = {1{`RANDOM}};
  way0Tag_81 = _RAND_209[20:0];
  _RAND_210 = {1{`RANDOM}};
  way0Tag_82 = _RAND_210[20:0];
  _RAND_211 = {1{`RANDOM}};
  way0Tag_83 = _RAND_211[20:0];
  _RAND_212 = {1{`RANDOM}};
  way0Tag_84 = _RAND_212[20:0];
  _RAND_213 = {1{`RANDOM}};
  way0Tag_85 = _RAND_213[20:0];
  _RAND_214 = {1{`RANDOM}};
  way0Tag_86 = _RAND_214[20:0];
  _RAND_215 = {1{`RANDOM}};
  way0Tag_87 = _RAND_215[20:0];
  _RAND_216 = {1{`RANDOM}};
  way0Tag_88 = _RAND_216[20:0];
  _RAND_217 = {1{`RANDOM}};
  way0Tag_89 = _RAND_217[20:0];
  _RAND_218 = {1{`RANDOM}};
  way0Tag_90 = _RAND_218[20:0];
  _RAND_219 = {1{`RANDOM}};
  way0Tag_91 = _RAND_219[20:0];
  _RAND_220 = {1{`RANDOM}};
  way0Tag_92 = _RAND_220[20:0];
  _RAND_221 = {1{`RANDOM}};
  way0Tag_93 = _RAND_221[20:0];
  _RAND_222 = {1{`RANDOM}};
  way0Tag_94 = _RAND_222[20:0];
  _RAND_223 = {1{`RANDOM}};
  way0Tag_95 = _RAND_223[20:0];
  _RAND_224 = {1{`RANDOM}};
  way0Tag_96 = _RAND_224[20:0];
  _RAND_225 = {1{`RANDOM}};
  way0Tag_97 = _RAND_225[20:0];
  _RAND_226 = {1{`RANDOM}};
  way0Tag_98 = _RAND_226[20:0];
  _RAND_227 = {1{`RANDOM}};
  way0Tag_99 = _RAND_227[20:0];
  _RAND_228 = {1{`RANDOM}};
  way0Tag_100 = _RAND_228[20:0];
  _RAND_229 = {1{`RANDOM}};
  way0Tag_101 = _RAND_229[20:0];
  _RAND_230 = {1{`RANDOM}};
  way0Tag_102 = _RAND_230[20:0];
  _RAND_231 = {1{`RANDOM}};
  way0Tag_103 = _RAND_231[20:0];
  _RAND_232 = {1{`RANDOM}};
  way0Tag_104 = _RAND_232[20:0];
  _RAND_233 = {1{`RANDOM}};
  way0Tag_105 = _RAND_233[20:0];
  _RAND_234 = {1{`RANDOM}};
  way0Tag_106 = _RAND_234[20:0];
  _RAND_235 = {1{`RANDOM}};
  way0Tag_107 = _RAND_235[20:0];
  _RAND_236 = {1{`RANDOM}};
  way0Tag_108 = _RAND_236[20:0];
  _RAND_237 = {1{`RANDOM}};
  way0Tag_109 = _RAND_237[20:0];
  _RAND_238 = {1{`RANDOM}};
  way0Tag_110 = _RAND_238[20:0];
  _RAND_239 = {1{`RANDOM}};
  way0Tag_111 = _RAND_239[20:0];
  _RAND_240 = {1{`RANDOM}};
  way0Tag_112 = _RAND_240[20:0];
  _RAND_241 = {1{`RANDOM}};
  way0Tag_113 = _RAND_241[20:0];
  _RAND_242 = {1{`RANDOM}};
  way0Tag_114 = _RAND_242[20:0];
  _RAND_243 = {1{`RANDOM}};
  way0Tag_115 = _RAND_243[20:0];
  _RAND_244 = {1{`RANDOM}};
  way0Tag_116 = _RAND_244[20:0];
  _RAND_245 = {1{`RANDOM}};
  way0Tag_117 = _RAND_245[20:0];
  _RAND_246 = {1{`RANDOM}};
  way0Tag_118 = _RAND_246[20:0];
  _RAND_247 = {1{`RANDOM}};
  way0Tag_119 = _RAND_247[20:0];
  _RAND_248 = {1{`RANDOM}};
  way0Tag_120 = _RAND_248[20:0];
  _RAND_249 = {1{`RANDOM}};
  way0Tag_121 = _RAND_249[20:0];
  _RAND_250 = {1{`RANDOM}};
  way0Tag_122 = _RAND_250[20:0];
  _RAND_251 = {1{`RANDOM}};
  way0Tag_123 = _RAND_251[20:0];
  _RAND_252 = {1{`RANDOM}};
  way0Tag_124 = _RAND_252[20:0];
  _RAND_253 = {1{`RANDOM}};
  way0Tag_125 = _RAND_253[20:0];
  _RAND_254 = {1{`RANDOM}};
  way0Tag_126 = _RAND_254[20:0];
  _RAND_255 = {1{`RANDOM}};
  way0Tag_127 = _RAND_255[20:0];
  _RAND_256 = {1{`RANDOM}};
  way0Age_0 = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  way0Age_1 = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  way0Age_2 = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  way0Age_3 = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  way0Age_4 = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  way0Age_5 = _RAND_261[0:0];
  _RAND_262 = {1{`RANDOM}};
  way0Age_6 = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  way0Age_7 = _RAND_263[0:0];
  _RAND_264 = {1{`RANDOM}};
  way0Age_8 = _RAND_264[0:0];
  _RAND_265 = {1{`RANDOM}};
  way0Age_9 = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  way0Age_10 = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  way0Age_11 = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  way0Age_12 = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  way0Age_13 = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  way0Age_14 = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  way0Age_15 = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  way0Age_16 = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  way0Age_17 = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  way0Age_18 = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  way0Age_19 = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  way0Age_20 = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  way0Age_21 = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  way0Age_22 = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  way0Age_23 = _RAND_279[0:0];
  _RAND_280 = {1{`RANDOM}};
  way0Age_24 = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  way0Age_25 = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  way0Age_26 = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  way0Age_27 = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  way0Age_28 = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  way0Age_29 = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  way0Age_30 = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  way0Age_31 = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  way0Age_32 = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  way0Age_33 = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  way0Age_34 = _RAND_290[0:0];
  _RAND_291 = {1{`RANDOM}};
  way0Age_35 = _RAND_291[0:0];
  _RAND_292 = {1{`RANDOM}};
  way0Age_36 = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  way0Age_37 = _RAND_293[0:0];
  _RAND_294 = {1{`RANDOM}};
  way0Age_38 = _RAND_294[0:0];
  _RAND_295 = {1{`RANDOM}};
  way0Age_39 = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  way0Age_40 = _RAND_296[0:0];
  _RAND_297 = {1{`RANDOM}};
  way0Age_41 = _RAND_297[0:0];
  _RAND_298 = {1{`RANDOM}};
  way0Age_42 = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  way0Age_43 = _RAND_299[0:0];
  _RAND_300 = {1{`RANDOM}};
  way0Age_44 = _RAND_300[0:0];
  _RAND_301 = {1{`RANDOM}};
  way0Age_45 = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  way0Age_46 = _RAND_302[0:0];
  _RAND_303 = {1{`RANDOM}};
  way0Age_47 = _RAND_303[0:0];
  _RAND_304 = {1{`RANDOM}};
  way0Age_48 = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  way0Age_49 = _RAND_305[0:0];
  _RAND_306 = {1{`RANDOM}};
  way0Age_50 = _RAND_306[0:0];
  _RAND_307 = {1{`RANDOM}};
  way0Age_51 = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  way0Age_52 = _RAND_308[0:0];
  _RAND_309 = {1{`RANDOM}};
  way0Age_53 = _RAND_309[0:0];
  _RAND_310 = {1{`RANDOM}};
  way0Age_54 = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  way0Age_55 = _RAND_311[0:0];
  _RAND_312 = {1{`RANDOM}};
  way0Age_56 = _RAND_312[0:0];
  _RAND_313 = {1{`RANDOM}};
  way0Age_57 = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  way0Age_58 = _RAND_314[0:0];
  _RAND_315 = {1{`RANDOM}};
  way0Age_59 = _RAND_315[0:0];
  _RAND_316 = {1{`RANDOM}};
  way0Age_60 = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  way0Age_61 = _RAND_317[0:0];
  _RAND_318 = {1{`RANDOM}};
  way0Age_62 = _RAND_318[0:0];
  _RAND_319 = {1{`RANDOM}};
  way0Age_63 = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  way0Age_64 = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  way0Age_65 = _RAND_321[0:0];
  _RAND_322 = {1{`RANDOM}};
  way0Age_66 = _RAND_322[0:0];
  _RAND_323 = {1{`RANDOM}};
  way0Age_67 = _RAND_323[0:0];
  _RAND_324 = {1{`RANDOM}};
  way0Age_68 = _RAND_324[0:0];
  _RAND_325 = {1{`RANDOM}};
  way0Age_69 = _RAND_325[0:0];
  _RAND_326 = {1{`RANDOM}};
  way0Age_70 = _RAND_326[0:0];
  _RAND_327 = {1{`RANDOM}};
  way0Age_71 = _RAND_327[0:0];
  _RAND_328 = {1{`RANDOM}};
  way0Age_72 = _RAND_328[0:0];
  _RAND_329 = {1{`RANDOM}};
  way0Age_73 = _RAND_329[0:0];
  _RAND_330 = {1{`RANDOM}};
  way0Age_74 = _RAND_330[0:0];
  _RAND_331 = {1{`RANDOM}};
  way0Age_75 = _RAND_331[0:0];
  _RAND_332 = {1{`RANDOM}};
  way0Age_76 = _RAND_332[0:0];
  _RAND_333 = {1{`RANDOM}};
  way0Age_77 = _RAND_333[0:0];
  _RAND_334 = {1{`RANDOM}};
  way0Age_78 = _RAND_334[0:0];
  _RAND_335 = {1{`RANDOM}};
  way0Age_79 = _RAND_335[0:0];
  _RAND_336 = {1{`RANDOM}};
  way0Age_80 = _RAND_336[0:0];
  _RAND_337 = {1{`RANDOM}};
  way0Age_81 = _RAND_337[0:0];
  _RAND_338 = {1{`RANDOM}};
  way0Age_82 = _RAND_338[0:0];
  _RAND_339 = {1{`RANDOM}};
  way0Age_83 = _RAND_339[0:0];
  _RAND_340 = {1{`RANDOM}};
  way0Age_84 = _RAND_340[0:0];
  _RAND_341 = {1{`RANDOM}};
  way0Age_85 = _RAND_341[0:0];
  _RAND_342 = {1{`RANDOM}};
  way0Age_86 = _RAND_342[0:0];
  _RAND_343 = {1{`RANDOM}};
  way0Age_87 = _RAND_343[0:0];
  _RAND_344 = {1{`RANDOM}};
  way0Age_88 = _RAND_344[0:0];
  _RAND_345 = {1{`RANDOM}};
  way0Age_89 = _RAND_345[0:0];
  _RAND_346 = {1{`RANDOM}};
  way0Age_90 = _RAND_346[0:0];
  _RAND_347 = {1{`RANDOM}};
  way0Age_91 = _RAND_347[0:0];
  _RAND_348 = {1{`RANDOM}};
  way0Age_92 = _RAND_348[0:0];
  _RAND_349 = {1{`RANDOM}};
  way0Age_93 = _RAND_349[0:0];
  _RAND_350 = {1{`RANDOM}};
  way0Age_94 = _RAND_350[0:0];
  _RAND_351 = {1{`RANDOM}};
  way0Age_95 = _RAND_351[0:0];
  _RAND_352 = {1{`RANDOM}};
  way0Age_96 = _RAND_352[0:0];
  _RAND_353 = {1{`RANDOM}};
  way0Age_97 = _RAND_353[0:0];
  _RAND_354 = {1{`RANDOM}};
  way0Age_98 = _RAND_354[0:0];
  _RAND_355 = {1{`RANDOM}};
  way0Age_99 = _RAND_355[0:0];
  _RAND_356 = {1{`RANDOM}};
  way0Age_100 = _RAND_356[0:0];
  _RAND_357 = {1{`RANDOM}};
  way0Age_101 = _RAND_357[0:0];
  _RAND_358 = {1{`RANDOM}};
  way0Age_102 = _RAND_358[0:0];
  _RAND_359 = {1{`RANDOM}};
  way0Age_103 = _RAND_359[0:0];
  _RAND_360 = {1{`RANDOM}};
  way0Age_104 = _RAND_360[0:0];
  _RAND_361 = {1{`RANDOM}};
  way0Age_105 = _RAND_361[0:0];
  _RAND_362 = {1{`RANDOM}};
  way0Age_106 = _RAND_362[0:0];
  _RAND_363 = {1{`RANDOM}};
  way0Age_107 = _RAND_363[0:0];
  _RAND_364 = {1{`RANDOM}};
  way0Age_108 = _RAND_364[0:0];
  _RAND_365 = {1{`RANDOM}};
  way0Age_109 = _RAND_365[0:0];
  _RAND_366 = {1{`RANDOM}};
  way0Age_110 = _RAND_366[0:0];
  _RAND_367 = {1{`RANDOM}};
  way0Age_111 = _RAND_367[0:0];
  _RAND_368 = {1{`RANDOM}};
  way0Age_112 = _RAND_368[0:0];
  _RAND_369 = {1{`RANDOM}};
  way0Age_113 = _RAND_369[0:0];
  _RAND_370 = {1{`RANDOM}};
  way0Age_114 = _RAND_370[0:0];
  _RAND_371 = {1{`RANDOM}};
  way0Age_115 = _RAND_371[0:0];
  _RAND_372 = {1{`RANDOM}};
  way0Age_116 = _RAND_372[0:0];
  _RAND_373 = {1{`RANDOM}};
  way0Age_117 = _RAND_373[0:0];
  _RAND_374 = {1{`RANDOM}};
  way0Age_118 = _RAND_374[0:0];
  _RAND_375 = {1{`RANDOM}};
  way0Age_119 = _RAND_375[0:0];
  _RAND_376 = {1{`RANDOM}};
  way0Age_120 = _RAND_376[0:0];
  _RAND_377 = {1{`RANDOM}};
  way0Age_121 = _RAND_377[0:0];
  _RAND_378 = {1{`RANDOM}};
  way0Age_122 = _RAND_378[0:0];
  _RAND_379 = {1{`RANDOM}};
  way0Age_123 = _RAND_379[0:0];
  _RAND_380 = {1{`RANDOM}};
  way0Age_124 = _RAND_380[0:0];
  _RAND_381 = {1{`RANDOM}};
  way0Age_125 = _RAND_381[0:0];
  _RAND_382 = {1{`RANDOM}};
  way0Age_126 = _RAND_382[0:0];
  _RAND_383 = {1{`RANDOM}};
  way0Age_127 = _RAND_383[0:0];
  _RAND_384 = {1{`RANDOM}};
  way0Dirty_0 = _RAND_384[0:0];
  _RAND_385 = {1{`RANDOM}};
  way0Dirty_1 = _RAND_385[0:0];
  _RAND_386 = {1{`RANDOM}};
  way0Dirty_2 = _RAND_386[0:0];
  _RAND_387 = {1{`RANDOM}};
  way0Dirty_3 = _RAND_387[0:0];
  _RAND_388 = {1{`RANDOM}};
  way0Dirty_4 = _RAND_388[0:0];
  _RAND_389 = {1{`RANDOM}};
  way0Dirty_5 = _RAND_389[0:0];
  _RAND_390 = {1{`RANDOM}};
  way0Dirty_6 = _RAND_390[0:0];
  _RAND_391 = {1{`RANDOM}};
  way0Dirty_7 = _RAND_391[0:0];
  _RAND_392 = {1{`RANDOM}};
  way0Dirty_8 = _RAND_392[0:0];
  _RAND_393 = {1{`RANDOM}};
  way0Dirty_9 = _RAND_393[0:0];
  _RAND_394 = {1{`RANDOM}};
  way0Dirty_10 = _RAND_394[0:0];
  _RAND_395 = {1{`RANDOM}};
  way0Dirty_11 = _RAND_395[0:0];
  _RAND_396 = {1{`RANDOM}};
  way0Dirty_12 = _RAND_396[0:0];
  _RAND_397 = {1{`RANDOM}};
  way0Dirty_13 = _RAND_397[0:0];
  _RAND_398 = {1{`RANDOM}};
  way0Dirty_14 = _RAND_398[0:0];
  _RAND_399 = {1{`RANDOM}};
  way0Dirty_15 = _RAND_399[0:0];
  _RAND_400 = {1{`RANDOM}};
  way0Dirty_16 = _RAND_400[0:0];
  _RAND_401 = {1{`RANDOM}};
  way0Dirty_17 = _RAND_401[0:0];
  _RAND_402 = {1{`RANDOM}};
  way0Dirty_18 = _RAND_402[0:0];
  _RAND_403 = {1{`RANDOM}};
  way0Dirty_19 = _RAND_403[0:0];
  _RAND_404 = {1{`RANDOM}};
  way0Dirty_20 = _RAND_404[0:0];
  _RAND_405 = {1{`RANDOM}};
  way0Dirty_21 = _RAND_405[0:0];
  _RAND_406 = {1{`RANDOM}};
  way0Dirty_22 = _RAND_406[0:0];
  _RAND_407 = {1{`RANDOM}};
  way0Dirty_23 = _RAND_407[0:0];
  _RAND_408 = {1{`RANDOM}};
  way0Dirty_24 = _RAND_408[0:0];
  _RAND_409 = {1{`RANDOM}};
  way0Dirty_25 = _RAND_409[0:0];
  _RAND_410 = {1{`RANDOM}};
  way0Dirty_26 = _RAND_410[0:0];
  _RAND_411 = {1{`RANDOM}};
  way0Dirty_27 = _RAND_411[0:0];
  _RAND_412 = {1{`RANDOM}};
  way0Dirty_28 = _RAND_412[0:0];
  _RAND_413 = {1{`RANDOM}};
  way0Dirty_29 = _RAND_413[0:0];
  _RAND_414 = {1{`RANDOM}};
  way0Dirty_30 = _RAND_414[0:0];
  _RAND_415 = {1{`RANDOM}};
  way0Dirty_31 = _RAND_415[0:0];
  _RAND_416 = {1{`RANDOM}};
  way0Dirty_32 = _RAND_416[0:0];
  _RAND_417 = {1{`RANDOM}};
  way0Dirty_33 = _RAND_417[0:0];
  _RAND_418 = {1{`RANDOM}};
  way0Dirty_34 = _RAND_418[0:0];
  _RAND_419 = {1{`RANDOM}};
  way0Dirty_35 = _RAND_419[0:0];
  _RAND_420 = {1{`RANDOM}};
  way0Dirty_36 = _RAND_420[0:0];
  _RAND_421 = {1{`RANDOM}};
  way0Dirty_37 = _RAND_421[0:0];
  _RAND_422 = {1{`RANDOM}};
  way0Dirty_38 = _RAND_422[0:0];
  _RAND_423 = {1{`RANDOM}};
  way0Dirty_39 = _RAND_423[0:0];
  _RAND_424 = {1{`RANDOM}};
  way0Dirty_40 = _RAND_424[0:0];
  _RAND_425 = {1{`RANDOM}};
  way0Dirty_41 = _RAND_425[0:0];
  _RAND_426 = {1{`RANDOM}};
  way0Dirty_42 = _RAND_426[0:0];
  _RAND_427 = {1{`RANDOM}};
  way0Dirty_43 = _RAND_427[0:0];
  _RAND_428 = {1{`RANDOM}};
  way0Dirty_44 = _RAND_428[0:0];
  _RAND_429 = {1{`RANDOM}};
  way0Dirty_45 = _RAND_429[0:0];
  _RAND_430 = {1{`RANDOM}};
  way0Dirty_46 = _RAND_430[0:0];
  _RAND_431 = {1{`RANDOM}};
  way0Dirty_47 = _RAND_431[0:0];
  _RAND_432 = {1{`RANDOM}};
  way0Dirty_48 = _RAND_432[0:0];
  _RAND_433 = {1{`RANDOM}};
  way0Dirty_49 = _RAND_433[0:0];
  _RAND_434 = {1{`RANDOM}};
  way0Dirty_50 = _RAND_434[0:0];
  _RAND_435 = {1{`RANDOM}};
  way0Dirty_51 = _RAND_435[0:0];
  _RAND_436 = {1{`RANDOM}};
  way0Dirty_52 = _RAND_436[0:0];
  _RAND_437 = {1{`RANDOM}};
  way0Dirty_53 = _RAND_437[0:0];
  _RAND_438 = {1{`RANDOM}};
  way0Dirty_54 = _RAND_438[0:0];
  _RAND_439 = {1{`RANDOM}};
  way0Dirty_55 = _RAND_439[0:0];
  _RAND_440 = {1{`RANDOM}};
  way0Dirty_56 = _RAND_440[0:0];
  _RAND_441 = {1{`RANDOM}};
  way0Dirty_57 = _RAND_441[0:0];
  _RAND_442 = {1{`RANDOM}};
  way0Dirty_58 = _RAND_442[0:0];
  _RAND_443 = {1{`RANDOM}};
  way0Dirty_59 = _RAND_443[0:0];
  _RAND_444 = {1{`RANDOM}};
  way0Dirty_60 = _RAND_444[0:0];
  _RAND_445 = {1{`RANDOM}};
  way0Dirty_61 = _RAND_445[0:0];
  _RAND_446 = {1{`RANDOM}};
  way0Dirty_62 = _RAND_446[0:0];
  _RAND_447 = {1{`RANDOM}};
  way0Dirty_63 = _RAND_447[0:0];
  _RAND_448 = {1{`RANDOM}};
  way0Dirty_64 = _RAND_448[0:0];
  _RAND_449 = {1{`RANDOM}};
  way0Dirty_65 = _RAND_449[0:0];
  _RAND_450 = {1{`RANDOM}};
  way0Dirty_66 = _RAND_450[0:0];
  _RAND_451 = {1{`RANDOM}};
  way0Dirty_67 = _RAND_451[0:0];
  _RAND_452 = {1{`RANDOM}};
  way0Dirty_68 = _RAND_452[0:0];
  _RAND_453 = {1{`RANDOM}};
  way0Dirty_69 = _RAND_453[0:0];
  _RAND_454 = {1{`RANDOM}};
  way0Dirty_70 = _RAND_454[0:0];
  _RAND_455 = {1{`RANDOM}};
  way0Dirty_71 = _RAND_455[0:0];
  _RAND_456 = {1{`RANDOM}};
  way0Dirty_72 = _RAND_456[0:0];
  _RAND_457 = {1{`RANDOM}};
  way0Dirty_73 = _RAND_457[0:0];
  _RAND_458 = {1{`RANDOM}};
  way0Dirty_74 = _RAND_458[0:0];
  _RAND_459 = {1{`RANDOM}};
  way0Dirty_75 = _RAND_459[0:0];
  _RAND_460 = {1{`RANDOM}};
  way0Dirty_76 = _RAND_460[0:0];
  _RAND_461 = {1{`RANDOM}};
  way0Dirty_77 = _RAND_461[0:0];
  _RAND_462 = {1{`RANDOM}};
  way0Dirty_78 = _RAND_462[0:0];
  _RAND_463 = {1{`RANDOM}};
  way0Dirty_79 = _RAND_463[0:0];
  _RAND_464 = {1{`RANDOM}};
  way0Dirty_80 = _RAND_464[0:0];
  _RAND_465 = {1{`RANDOM}};
  way0Dirty_81 = _RAND_465[0:0];
  _RAND_466 = {1{`RANDOM}};
  way0Dirty_82 = _RAND_466[0:0];
  _RAND_467 = {1{`RANDOM}};
  way0Dirty_83 = _RAND_467[0:0];
  _RAND_468 = {1{`RANDOM}};
  way0Dirty_84 = _RAND_468[0:0];
  _RAND_469 = {1{`RANDOM}};
  way0Dirty_85 = _RAND_469[0:0];
  _RAND_470 = {1{`RANDOM}};
  way0Dirty_86 = _RAND_470[0:0];
  _RAND_471 = {1{`RANDOM}};
  way0Dirty_87 = _RAND_471[0:0];
  _RAND_472 = {1{`RANDOM}};
  way0Dirty_88 = _RAND_472[0:0];
  _RAND_473 = {1{`RANDOM}};
  way0Dirty_89 = _RAND_473[0:0];
  _RAND_474 = {1{`RANDOM}};
  way0Dirty_90 = _RAND_474[0:0];
  _RAND_475 = {1{`RANDOM}};
  way0Dirty_91 = _RAND_475[0:0];
  _RAND_476 = {1{`RANDOM}};
  way0Dirty_92 = _RAND_476[0:0];
  _RAND_477 = {1{`RANDOM}};
  way0Dirty_93 = _RAND_477[0:0];
  _RAND_478 = {1{`RANDOM}};
  way0Dirty_94 = _RAND_478[0:0];
  _RAND_479 = {1{`RANDOM}};
  way0Dirty_95 = _RAND_479[0:0];
  _RAND_480 = {1{`RANDOM}};
  way0Dirty_96 = _RAND_480[0:0];
  _RAND_481 = {1{`RANDOM}};
  way0Dirty_97 = _RAND_481[0:0];
  _RAND_482 = {1{`RANDOM}};
  way0Dirty_98 = _RAND_482[0:0];
  _RAND_483 = {1{`RANDOM}};
  way0Dirty_99 = _RAND_483[0:0];
  _RAND_484 = {1{`RANDOM}};
  way0Dirty_100 = _RAND_484[0:0];
  _RAND_485 = {1{`RANDOM}};
  way0Dirty_101 = _RAND_485[0:0];
  _RAND_486 = {1{`RANDOM}};
  way0Dirty_102 = _RAND_486[0:0];
  _RAND_487 = {1{`RANDOM}};
  way0Dirty_103 = _RAND_487[0:0];
  _RAND_488 = {1{`RANDOM}};
  way0Dirty_104 = _RAND_488[0:0];
  _RAND_489 = {1{`RANDOM}};
  way0Dirty_105 = _RAND_489[0:0];
  _RAND_490 = {1{`RANDOM}};
  way0Dirty_106 = _RAND_490[0:0];
  _RAND_491 = {1{`RANDOM}};
  way0Dirty_107 = _RAND_491[0:0];
  _RAND_492 = {1{`RANDOM}};
  way0Dirty_108 = _RAND_492[0:0];
  _RAND_493 = {1{`RANDOM}};
  way0Dirty_109 = _RAND_493[0:0];
  _RAND_494 = {1{`RANDOM}};
  way0Dirty_110 = _RAND_494[0:0];
  _RAND_495 = {1{`RANDOM}};
  way0Dirty_111 = _RAND_495[0:0];
  _RAND_496 = {1{`RANDOM}};
  way0Dirty_112 = _RAND_496[0:0];
  _RAND_497 = {1{`RANDOM}};
  way0Dirty_113 = _RAND_497[0:0];
  _RAND_498 = {1{`RANDOM}};
  way0Dirty_114 = _RAND_498[0:0];
  _RAND_499 = {1{`RANDOM}};
  way0Dirty_115 = _RAND_499[0:0];
  _RAND_500 = {1{`RANDOM}};
  way0Dirty_116 = _RAND_500[0:0];
  _RAND_501 = {1{`RANDOM}};
  way0Dirty_117 = _RAND_501[0:0];
  _RAND_502 = {1{`RANDOM}};
  way0Dirty_118 = _RAND_502[0:0];
  _RAND_503 = {1{`RANDOM}};
  way0Dirty_119 = _RAND_503[0:0];
  _RAND_504 = {1{`RANDOM}};
  way0Dirty_120 = _RAND_504[0:0];
  _RAND_505 = {1{`RANDOM}};
  way0Dirty_121 = _RAND_505[0:0];
  _RAND_506 = {1{`RANDOM}};
  way0Dirty_122 = _RAND_506[0:0];
  _RAND_507 = {1{`RANDOM}};
  way0Dirty_123 = _RAND_507[0:0];
  _RAND_508 = {1{`RANDOM}};
  way0Dirty_124 = _RAND_508[0:0];
  _RAND_509 = {1{`RANDOM}};
  way0Dirty_125 = _RAND_509[0:0];
  _RAND_510 = {1{`RANDOM}};
  way0Dirty_126 = _RAND_510[0:0];
  _RAND_511 = {1{`RANDOM}};
  way0Dirty_127 = _RAND_511[0:0];
  _RAND_512 = {1{`RANDOM}};
  way1V_0 = _RAND_512[0:0];
  _RAND_513 = {1{`RANDOM}};
  way1V_1 = _RAND_513[0:0];
  _RAND_514 = {1{`RANDOM}};
  way1V_2 = _RAND_514[0:0];
  _RAND_515 = {1{`RANDOM}};
  way1V_3 = _RAND_515[0:0];
  _RAND_516 = {1{`RANDOM}};
  way1V_4 = _RAND_516[0:0];
  _RAND_517 = {1{`RANDOM}};
  way1V_5 = _RAND_517[0:0];
  _RAND_518 = {1{`RANDOM}};
  way1V_6 = _RAND_518[0:0];
  _RAND_519 = {1{`RANDOM}};
  way1V_7 = _RAND_519[0:0];
  _RAND_520 = {1{`RANDOM}};
  way1V_8 = _RAND_520[0:0];
  _RAND_521 = {1{`RANDOM}};
  way1V_9 = _RAND_521[0:0];
  _RAND_522 = {1{`RANDOM}};
  way1V_10 = _RAND_522[0:0];
  _RAND_523 = {1{`RANDOM}};
  way1V_11 = _RAND_523[0:0];
  _RAND_524 = {1{`RANDOM}};
  way1V_12 = _RAND_524[0:0];
  _RAND_525 = {1{`RANDOM}};
  way1V_13 = _RAND_525[0:0];
  _RAND_526 = {1{`RANDOM}};
  way1V_14 = _RAND_526[0:0];
  _RAND_527 = {1{`RANDOM}};
  way1V_15 = _RAND_527[0:0];
  _RAND_528 = {1{`RANDOM}};
  way1V_16 = _RAND_528[0:0];
  _RAND_529 = {1{`RANDOM}};
  way1V_17 = _RAND_529[0:0];
  _RAND_530 = {1{`RANDOM}};
  way1V_18 = _RAND_530[0:0];
  _RAND_531 = {1{`RANDOM}};
  way1V_19 = _RAND_531[0:0];
  _RAND_532 = {1{`RANDOM}};
  way1V_20 = _RAND_532[0:0];
  _RAND_533 = {1{`RANDOM}};
  way1V_21 = _RAND_533[0:0];
  _RAND_534 = {1{`RANDOM}};
  way1V_22 = _RAND_534[0:0];
  _RAND_535 = {1{`RANDOM}};
  way1V_23 = _RAND_535[0:0];
  _RAND_536 = {1{`RANDOM}};
  way1V_24 = _RAND_536[0:0];
  _RAND_537 = {1{`RANDOM}};
  way1V_25 = _RAND_537[0:0];
  _RAND_538 = {1{`RANDOM}};
  way1V_26 = _RAND_538[0:0];
  _RAND_539 = {1{`RANDOM}};
  way1V_27 = _RAND_539[0:0];
  _RAND_540 = {1{`RANDOM}};
  way1V_28 = _RAND_540[0:0];
  _RAND_541 = {1{`RANDOM}};
  way1V_29 = _RAND_541[0:0];
  _RAND_542 = {1{`RANDOM}};
  way1V_30 = _RAND_542[0:0];
  _RAND_543 = {1{`RANDOM}};
  way1V_31 = _RAND_543[0:0];
  _RAND_544 = {1{`RANDOM}};
  way1V_32 = _RAND_544[0:0];
  _RAND_545 = {1{`RANDOM}};
  way1V_33 = _RAND_545[0:0];
  _RAND_546 = {1{`RANDOM}};
  way1V_34 = _RAND_546[0:0];
  _RAND_547 = {1{`RANDOM}};
  way1V_35 = _RAND_547[0:0];
  _RAND_548 = {1{`RANDOM}};
  way1V_36 = _RAND_548[0:0];
  _RAND_549 = {1{`RANDOM}};
  way1V_37 = _RAND_549[0:0];
  _RAND_550 = {1{`RANDOM}};
  way1V_38 = _RAND_550[0:0];
  _RAND_551 = {1{`RANDOM}};
  way1V_39 = _RAND_551[0:0];
  _RAND_552 = {1{`RANDOM}};
  way1V_40 = _RAND_552[0:0];
  _RAND_553 = {1{`RANDOM}};
  way1V_41 = _RAND_553[0:0];
  _RAND_554 = {1{`RANDOM}};
  way1V_42 = _RAND_554[0:0];
  _RAND_555 = {1{`RANDOM}};
  way1V_43 = _RAND_555[0:0];
  _RAND_556 = {1{`RANDOM}};
  way1V_44 = _RAND_556[0:0];
  _RAND_557 = {1{`RANDOM}};
  way1V_45 = _RAND_557[0:0];
  _RAND_558 = {1{`RANDOM}};
  way1V_46 = _RAND_558[0:0];
  _RAND_559 = {1{`RANDOM}};
  way1V_47 = _RAND_559[0:0];
  _RAND_560 = {1{`RANDOM}};
  way1V_48 = _RAND_560[0:0];
  _RAND_561 = {1{`RANDOM}};
  way1V_49 = _RAND_561[0:0];
  _RAND_562 = {1{`RANDOM}};
  way1V_50 = _RAND_562[0:0];
  _RAND_563 = {1{`RANDOM}};
  way1V_51 = _RAND_563[0:0];
  _RAND_564 = {1{`RANDOM}};
  way1V_52 = _RAND_564[0:0];
  _RAND_565 = {1{`RANDOM}};
  way1V_53 = _RAND_565[0:0];
  _RAND_566 = {1{`RANDOM}};
  way1V_54 = _RAND_566[0:0];
  _RAND_567 = {1{`RANDOM}};
  way1V_55 = _RAND_567[0:0];
  _RAND_568 = {1{`RANDOM}};
  way1V_56 = _RAND_568[0:0];
  _RAND_569 = {1{`RANDOM}};
  way1V_57 = _RAND_569[0:0];
  _RAND_570 = {1{`RANDOM}};
  way1V_58 = _RAND_570[0:0];
  _RAND_571 = {1{`RANDOM}};
  way1V_59 = _RAND_571[0:0];
  _RAND_572 = {1{`RANDOM}};
  way1V_60 = _RAND_572[0:0];
  _RAND_573 = {1{`RANDOM}};
  way1V_61 = _RAND_573[0:0];
  _RAND_574 = {1{`RANDOM}};
  way1V_62 = _RAND_574[0:0];
  _RAND_575 = {1{`RANDOM}};
  way1V_63 = _RAND_575[0:0];
  _RAND_576 = {1{`RANDOM}};
  way1V_64 = _RAND_576[0:0];
  _RAND_577 = {1{`RANDOM}};
  way1V_65 = _RAND_577[0:0];
  _RAND_578 = {1{`RANDOM}};
  way1V_66 = _RAND_578[0:0];
  _RAND_579 = {1{`RANDOM}};
  way1V_67 = _RAND_579[0:0];
  _RAND_580 = {1{`RANDOM}};
  way1V_68 = _RAND_580[0:0];
  _RAND_581 = {1{`RANDOM}};
  way1V_69 = _RAND_581[0:0];
  _RAND_582 = {1{`RANDOM}};
  way1V_70 = _RAND_582[0:0];
  _RAND_583 = {1{`RANDOM}};
  way1V_71 = _RAND_583[0:0];
  _RAND_584 = {1{`RANDOM}};
  way1V_72 = _RAND_584[0:0];
  _RAND_585 = {1{`RANDOM}};
  way1V_73 = _RAND_585[0:0];
  _RAND_586 = {1{`RANDOM}};
  way1V_74 = _RAND_586[0:0];
  _RAND_587 = {1{`RANDOM}};
  way1V_75 = _RAND_587[0:0];
  _RAND_588 = {1{`RANDOM}};
  way1V_76 = _RAND_588[0:0];
  _RAND_589 = {1{`RANDOM}};
  way1V_77 = _RAND_589[0:0];
  _RAND_590 = {1{`RANDOM}};
  way1V_78 = _RAND_590[0:0];
  _RAND_591 = {1{`RANDOM}};
  way1V_79 = _RAND_591[0:0];
  _RAND_592 = {1{`RANDOM}};
  way1V_80 = _RAND_592[0:0];
  _RAND_593 = {1{`RANDOM}};
  way1V_81 = _RAND_593[0:0];
  _RAND_594 = {1{`RANDOM}};
  way1V_82 = _RAND_594[0:0];
  _RAND_595 = {1{`RANDOM}};
  way1V_83 = _RAND_595[0:0];
  _RAND_596 = {1{`RANDOM}};
  way1V_84 = _RAND_596[0:0];
  _RAND_597 = {1{`RANDOM}};
  way1V_85 = _RAND_597[0:0];
  _RAND_598 = {1{`RANDOM}};
  way1V_86 = _RAND_598[0:0];
  _RAND_599 = {1{`RANDOM}};
  way1V_87 = _RAND_599[0:0];
  _RAND_600 = {1{`RANDOM}};
  way1V_88 = _RAND_600[0:0];
  _RAND_601 = {1{`RANDOM}};
  way1V_89 = _RAND_601[0:0];
  _RAND_602 = {1{`RANDOM}};
  way1V_90 = _RAND_602[0:0];
  _RAND_603 = {1{`RANDOM}};
  way1V_91 = _RAND_603[0:0];
  _RAND_604 = {1{`RANDOM}};
  way1V_92 = _RAND_604[0:0];
  _RAND_605 = {1{`RANDOM}};
  way1V_93 = _RAND_605[0:0];
  _RAND_606 = {1{`RANDOM}};
  way1V_94 = _RAND_606[0:0];
  _RAND_607 = {1{`RANDOM}};
  way1V_95 = _RAND_607[0:0];
  _RAND_608 = {1{`RANDOM}};
  way1V_96 = _RAND_608[0:0];
  _RAND_609 = {1{`RANDOM}};
  way1V_97 = _RAND_609[0:0];
  _RAND_610 = {1{`RANDOM}};
  way1V_98 = _RAND_610[0:0];
  _RAND_611 = {1{`RANDOM}};
  way1V_99 = _RAND_611[0:0];
  _RAND_612 = {1{`RANDOM}};
  way1V_100 = _RAND_612[0:0];
  _RAND_613 = {1{`RANDOM}};
  way1V_101 = _RAND_613[0:0];
  _RAND_614 = {1{`RANDOM}};
  way1V_102 = _RAND_614[0:0];
  _RAND_615 = {1{`RANDOM}};
  way1V_103 = _RAND_615[0:0];
  _RAND_616 = {1{`RANDOM}};
  way1V_104 = _RAND_616[0:0];
  _RAND_617 = {1{`RANDOM}};
  way1V_105 = _RAND_617[0:0];
  _RAND_618 = {1{`RANDOM}};
  way1V_106 = _RAND_618[0:0];
  _RAND_619 = {1{`RANDOM}};
  way1V_107 = _RAND_619[0:0];
  _RAND_620 = {1{`RANDOM}};
  way1V_108 = _RAND_620[0:0];
  _RAND_621 = {1{`RANDOM}};
  way1V_109 = _RAND_621[0:0];
  _RAND_622 = {1{`RANDOM}};
  way1V_110 = _RAND_622[0:0];
  _RAND_623 = {1{`RANDOM}};
  way1V_111 = _RAND_623[0:0];
  _RAND_624 = {1{`RANDOM}};
  way1V_112 = _RAND_624[0:0];
  _RAND_625 = {1{`RANDOM}};
  way1V_113 = _RAND_625[0:0];
  _RAND_626 = {1{`RANDOM}};
  way1V_114 = _RAND_626[0:0];
  _RAND_627 = {1{`RANDOM}};
  way1V_115 = _RAND_627[0:0];
  _RAND_628 = {1{`RANDOM}};
  way1V_116 = _RAND_628[0:0];
  _RAND_629 = {1{`RANDOM}};
  way1V_117 = _RAND_629[0:0];
  _RAND_630 = {1{`RANDOM}};
  way1V_118 = _RAND_630[0:0];
  _RAND_631 = {1{`RANDOM}};
  way1V_119 = _RAND_631[0:0];
  _RAND_632 = {1{`RANDOM}};
  way1V_120 = _RAND_632[0:0];
  _RAND_633 = {1{`RANDOM}};
  way1V_121 = _RAND_633[0:0];
  _RAND_634 = {1{`RANDOM}};
  way1V_122 = _RAND_634[0:0];
  _RAND_635 = {1{`RANDOM}};
  way1V_123 = _RAND_635[0:0];
  _RAND_636 = {1{`RANDOM}};
  way1V_124 = _RAND_636[0:0];
  _RAND_637 = {1{`RANDOM}};
  way1V_125 = _RAND_637[0:0];
  _RAND_638 = {1{`RANDOM}};
  way1V_126 = _RAND_638[0:0];
  _RAND_639 = {1{`RANDOM}};
  way1V_127 = _RAND_639[0:0];
  _RAND_640 = {1{`RANDOM}};
  way1Tag_0 = _RAND_640[20:0];
  _RAND_641 = {1{`RANDOM}};
  way1Tag_1 = _RAND_641[20:0];
  _RAND_642 = {1{`RANDOM}};
  way1Tag_2 = _RAND_642[20:0];
  _RAND_643 = {1{`RANDOM}};
  way1Tag_3 = _RAND_643[20:0];
  _RAND_644 = {1{`RANDOM}};
  way1Tag_4 = _RAND_644[20:0];
  _RAND_645 = {1{`RANDOM}};
  way1Tag_5 = _RAND_645[20:0];
  _RAND_646 = {1{`RANDOM}};
  way1Tag_6 = _RAND_646[20:0];
  _RAND_647 = {1{`RANDOM}};
  way1Tag_7 = _RAND_647[20:0];
  _RAND_648 = {1{`RANDOM}};
  way1Tag_8 = _RAND_648[20:0];
  _RAND_649 = {1{`RANDOM}};
  way1Tag_9 = _RAND_649[20:0];
  _RAND_650 = {1{`RANDOM}};
  way1Tag_10 = _RAND_650[20:0];
  _RAND_651 = {1{`RANDOM}};
  way1Tag_11 = _RAND_651[20:0];
  _RAND_652 = {1{`RANDOM}};
  way1Tag_12 = _RAND_652[20:0];
  _RAND_653 = {1{`RANDOM}};
  way1Tag_13 = _RAND_653[20:0];
  _RAND_654 = {1{`RANDOM}};
  way1Tag_14 = _RAND_654[20:0];
  _RAND_655 = {1{`RANDOM}};
  way1Tag_15 = _RAND_655[20:0];
  _RAND_656 = {1{`RANDOM}};
  way1Tag_16 = _RAND_656[20:0];
  _RAND_657 = {1{`RANDOM}};
  way1Tag_17 = _RAND_657[20:0];
  _RAND_658 = {1{`RANDOM}};
  way1Tag_18 = _RAND_658[20:0];
  _RAND_659 = {1{`RANDOM}};
  way1Tag_19 = _RAND_659[20:0];
  _RAND_660 = {1{`RANDOM}};
  way1Tag_20 = _RAND_660[20:0];
  _RAND_661 = {1{`RANDOM}};
  way1Tag_21 = _RAND_661[20:0];
  _RAND_662 = {1{`RANDOM}};
  way1Tag_22 = _RAND_662[20:0];
  _RAND_663 = {1{`RANDOM}};
  way1Tag_23 = _RAND_663[20:0];
  _RAND_664 = {1{`RANDOM}};
  way1Tag_24 = _RAND_664[20:0];
  _RAND_665 = {1{`RANDOM}};
  way1Tag_25 = _RAND_665[20:0];
  _RAND_666 = {1{`RANDOM}};
  way1Tag_26 = _RAND_666[20:0];
  _RAND_667 = {1{`RANDOM}};
  way1Tag_27 = _RAND_667[20:0];
  _RAND_668 = {1{`RANDOM}};
  way1Tag_28 = _RAND_668[20:0];
  _RAND_669 = {1{`RANDOM}};
  way1Tag_29 = _RAND_669[20:0];
  _RAND_670 = {1{`RANDOM}};
  way1Tag_30 = _RAND_670[20:0];
  _RAND_671 = {1{`RANDOM}};
  way1Tag_31 = _RAND_671[20:0];
  _RAND_672 = {1{`RANDOM}};
  way1Tag_32 = _RAND_672[20:0];
  _RAND_673 = {1{`RANDOM}};
  way1Tag_33 = _RAND_673[20:0];
  _RAND_674 = {1{`RANDOM}};
  way1Tag_34 = _RAND_674[20:0];
  _RAND_675 = {1{`RANDOM}};
  way1Tag_35 = _RAND_675[20:0];
  _RAND_676 = {1{`RANDOM}};
  way1Tag_36 = _RAND_676[20:0];
  _RAND_677 = {1{`RANDOM}};
  way1Tag_37 = _RAND_677[20:0];
  _RAND_678 = {1{`RANDOM}};
  way1Tag_38 = _RAND_678[20:0];
  _RAND_679 = {1{`RANDOM}};
  way1Tag_39 = _RAND_679[20:0];
  _RAND_680 = {1{`RANDOM}};
  way1Tag_40 = _RAND_680[20:0];
  _RAND_681 = {1{`RANDOM}};
  way1Tag_41 = _RAND_681[20:0];
  _RAND_682 = {1{`RANDOM}};
  way1Tag_42 = _RAND_682[20:0];
  _RAND_683 = {1{`RANDOM}};
  way1Tag_43 = _RAND_683[20:0];
  _RAND_684 = {1{`RANDOM}};
  way1Tag_44 = _RAND_684[20:0];
  _RAND_685 = {1{`RANDOM}};
  way1Tag_45 = _RAND_685[20:0];
  _RAND_686 = {1{`RANDOM}};
  way1Tag_46 = _RAND_686[20:0];
  _RAND_687 = {1{`RANDOM}};
  way1Tag_47 = _RAND_687[20:0];
  _RAND_688 = {1{`RANDOM}};
  way1Tag_48 = _RAND_688[20:0];
  _RAND_689 = {1{`RANDOM}};
  way1Tag_49 = _RAND_689[20:0];
  _RAND_690 = {1{`RANDOM}};
  way1Tag_50 = _RAND_690[20:0];
  _RAND_691 = {1{`RANDOM}};
  way1Tag_51 = _RAND_691[20:0];
  _RAND_692 = {1{`RANDOM}};
  way1Tag_52 = _RAND_692[20:0];
  _RAND_693 = {1{`RANDOM}};
  way1Tag_53 = _RAND_693[20:0];
  _RAND_694 = {1{`RANDOM}};
  way1Tag_54 = _RAND_694[20:0];
  _RAND_695 = {1{`RANDOM}};
  way1Tag_55 = _RAND_695[20:0];
  _RAND_696 = {1{`RANDOM}};
  way1Tag_56 = _RAND_696[20:0];
  _RAND_697 = {1{`RANDOM}};
  way1Tag_57 = _RAND_697[20:0];
  _RAND_698 = {1{`RANDOM}};
  way1Tag_58 = _RAND_698[20:0];
  _RAND_699 = {1{`RANDOM}};
  way1Tag_59 = _RAND_699[20:0];
  _RAND_700 = {1{`RANDOM}};
  way1Tag_60 = _RAND_700[20:0];
  _RAND_701 = {1{`RANDOM}};
  way1Tag_61 = _RAND_701[20:0];
  _RAND_702 = {1{`RANDOM}};
  way1Tag_62 = _RAND_702[20:0];
  _RAND_703 = {1{`RANDOM}};
  way1Tag_63 = _RAND_703[20:0];
  _RAND_704 = {1{`RANDOM}};
  way1Tag_64 = _RAND_704[20:0];
  _RAND_705 = {1{`RANDOM}};
  way1Tag_65 = _RAND_705[20:0];
  _RAND_706 = {1{`RANDOM}};
  way1Tag_66 = _RAND_706[20:0];
  _RAND_707 = {1{`RANDOM}};
  way1Tag_67 = _RAND_707[20:0];
  _RAND_708 = {1{`RANDOM}};
  way1Tag_68 = _RAND_708[20:0];
  _RAND_709 = {1{`RANDOM}};
  way1Tag_69 = _RAND_709[20:0];
  _RAND_710 = {1{`RANDOM}};
  way1Tag_70 = _RAND_710[20:0];
  _RAND_711 = {1{`RANDOM}};
  way1Tag_71 = _RAND_711[20:0];
  _RAND_712 = {1{`RANDOM}};
  way1Tag_72 = _RAND_712[20:0];
  _RAND_713 = {1{`RANDOM}};
  way1Tag_73 = _RAND_713[20:0];
  _RAND_714 = {1{`RANDOM}};
  way1Tag_74 = _RAND_714[20:0];
  _RAND_715 = {1{`RANDOM}};
  way1Tag_75 = _RAND_715[20:0];
  _RAND_716 = {1{`RANDOM}};
  way1Tag_76 = _RAND_716[20:0];
  _RAND_717 = {1{`RANDOM}};
  way1Tag_77 = _RAND_717[20:0];
  _RAND_718 = {1{`RANDOM}};
  way1Tag_78 = _RAND_718[20:0];
  _RAND_719 = {1{`RANDOM}};
  way1Tag_79 = _RAND_719[20:0];
  _RAND_720 = {1{`RANDOM}};
  way1Tag_80 = _RAND_720[20:0];
  _RAND_721 = {1{`RANDOM}};
  way1Tag_81 = _RAND_721[20:0];
  _RAND_722 = {1{`RANDOM}};
  way1Tag_82 = _RAND_722[20:0];
  _RAND_723 = {1{`RANDOM}};
  way1Tag_83 = _RAND_723[20:0];
  _RAND_724 = {1{`RANDOM}};
  way1Tag_84 = _RAND_724[20:0];
  _RAND_725 = {1{`RANDOM}};
  way1Tag_85 = _RAND_725[20:0];
  _RAND_726 = {1{`RANDOM}};
  way1Tag_86 = _RAND_726[20:0];
  _RAND_727 = {1{`RANDOM}};
  way1Tag_87 = _RAND_727[20:0];
  _RAND_728 = {1{`RANDOM}};
  way1Tag_88 = _RAND_728[20:0];
  _RAND_729 = {1{`RANDOM}};
  way1Tag_89 = _RAND_729[20:0];
  _RAND_730 = {1{`RANDOM}};
  way1Tag_90 = _RAND_730[20:0];
  _RAND_731 = {1{`RANDOM}};
  way1Tag_91 = _RAND_731[20:0];
  _RAND_732 = {1{`RANDOM}};
  way1Tag_92 = _RAND_732[20:0];
  _RAND_733 = {1{`RANDOM}};
  way1Tag_93 = _RAND_733[20:0];
  _RAND_734 = {1{`RANDOM}};
  way1Tag_94 = _RAND_734[20:0];
  _RAND_735 = {1{`RANDOM}};
  way1Tag_95 = _RAND_735[20:0];
  _RAND_736 = {1{`RANDOM}};
  way1Tag_96 = _RAND_736[20:0];
  _RAND_737 = {1{`RANDOM}};
  way1Tag_97 = _RAND_737[20:0];
  _RAND_738 = {1{`RANDOM}};
  way1Tag_98 = _RAND_738[20:0];
  _RAND_739 = {1{`RANDOM}};
  way1Tag_99 = _RAND_739[20:0];
  _RAND_740 = {1{`RANDOM}};
  way1Tag_100 = _RAND_740[20:0];
  _RAND_741 = {1{`RANDOM}};
  way1Tag_101 = _RAND_741[20:0];
  _RAND_742 = {1{`RANDOM}};
  way1Tag_102 = _RAND_742[20:0];
  _RAND_743 = {1{`RANDOM}};
  way1Tag_103 = _RAND_743[20:0];
  _RAND_744 = {1{`RANDOM}};
  way1Tag_104 = _RAND_744[20:0];
  _RAND_745 = {1{`RANDOM}};
  way1Tag_105 = _RAND_745[20:0];
  _RAND_746 = {1{`RANDOM}};
  way1Tag_106 = _RAND_746[20:0];
  _RAND_747 = {1{`RANDOM}};
  way1Tag_107 = _RAND_747[20:0];
  _RAND_748 = {1{`RANDOM}};
  way1Tag_108 = _RAND_748[20:0];
  _RAND_749 = {1{`RANDOM}};
  way1Tag_109 = _RAND_749[20:0];
  _RAND_750 = {1{`RANDOM}};
  way1Tag_110 = _RAND_750[20:0];
  _RAND_751 = {1{`RANDOM}};
  way1Tag_111 = _RAND_751[20:0];
  _RAND_752 = {1{`RANDOM}};
  way1Tag_112 = _RAND_752[20:0];
  _RAND_753 = {1{`RANDOM}};
  way1Tag_113 = _RAND_753[20:0];
  _RAND_754 = {1{`RANDOM}};
  way1Tag_114 = _RAND_754[20:0];
  _RAND_755 = {1{`RANDOM}};
  way1Tag_115 = _RAND_755[20:0];
  _RAND_756 = {1{`RANDOM}};
  way1Tag_116 = _RAND_756[20:0];
  _RAND_757 = {1{`RANDOM}};
  way1Tag_117 = _RAND_757[20:0];
  _RAND_758 = {1{`RANDOM}};
  way1Tag_118 = _RAND_758[20:0];
  _RAND_759 = {1{`RANDOM}};
  way1Tag_119 = _RAND_759[20:0];
  _RAND_760 = {1{`RANDOM}};
  way1Tag_120 = _RAND_760[20:0];
  _RAND_761 = {1{`RANDOM}};
  way1Tag_121 = _RAND_761[20:0];
  _RAND_762 = {1{`RANDOM}};
  way1Tag_122 = _RAND_762[20:0];
  _RAND_763 = {1{`RANDOM}};
  way1Tag_123 = _RAND_763[20:0];
  _RAND_764 = {1{`RANDOM}};
  way1Tag_124 = _RAND_764[20:0];
  _RAND_765 = {1{`RANDOM}};
  way1Tag_125 = _RAND_765[20:0];
  _RAND_766 = {1{`RANDOM}};
  way1Tag_126 = _RAND_766[20:0];
  _RAND_767 = {1{`RANDOM}};
  way1Tag_127 = _RAND_767[20:0];
  _RAND_768 = {1{`RANDOM}};
  way1Dirty_0 = _RAND_768[0:0];
  _RAND_769 = {1{`RANDOM}};
  way1Dirty_1 = _RAND_769[0:0];
  _RAND_770 = {1{`RANDOM}};
  way1Dirty_2 = _RAND_770[0:0];
  _RAND_771 = {1{`RANDOM}};
  way1Dirty_3 = _RAND_771[0:0];
  _RAND_772 = {1{`RANDOM}};
  way1Dirty_4 = _RAND_772[0:0];
  _RAND_773 = {1{`RANDOM}};
  way1Dirty_5 = _RAND_773[0:0];
  _RAND_774 = {1{`RANDOM}};
  way1Dirty_6 = _RAND_774[0:0];
  _RAND_775 = {1{`RANDOM}};
  way1Dirty_7 = _RAND_775[0:0];
  _RAND_776 = {1{`RANDOM}};
  way1Dirty_8 = _RAND_776[0:0];
  _RAND_777 = {1{`RANDOM}};
  way1Dirty_9 = _RAND_777[0:0];
  _RAND_778 = {1{`RANDOM}};
  way1Dirty_10 = _RAND_778[0:0];
  _RAND_779 = {1{`RANDOM}};
  way1Dirty_11 = _RAND_779[0:0];
  _RAND_780 = {1{`RANDOM}};
  way1Dirty_12 = _RAND_780[0:0];
  _RAND_781 = {1{`RANDOM}};
  way1Dirty_13 = _RAND_781[0:0];
  _RAND_782 = {1{`RANDOM}};
  way1Dirty_14 = _RAND_782[0:0];
  _RAND_783 = {1{`RANDOM}};
  way1Dirty_15 = _RAND_783[0:0];
  _RAND_784 = {1{`RANDOM}};
  way1Dirty_16 = _RAND_784[0:0];
  _RAND_785 = {1{`RANDOM}};
  way1Dirty_17 = _RAND_785[0:0];
  _RAND_786 = {1{`RANDOM}};
  way1Dirty_18 = _RAND_786[0:0];
  _RAND_787 = {1{`RANDOM}};
  way1Dirty_19 = _RAND_787[0:0];
  _RAND_788 = {1{`RANDOM}};
  way1Dirty_20 = _RAND_788[0:0];
  _RAND_789 = {1{`RANDOM}};
  way1Dirty_21 = _RAND_789[0:0];
  _RAND_790 = {1{`RANDOM}};
  way1Dirty_22 = _RAND_790[0:0];
  _RAND_791 = {1{`RANDOM}};
  way1Dirty_23 = _RAND_791[0:0];
  _RAND_792 = {1{`RANDOM}};
  way1Dirty_24 = _RAND_792[0:0];
  _RAND_793 = {1{`RANDOM}};
  way1Dirty_25 = _RAND_793[0:0];
  _RAND_794 = {1{`RANDOM}};
  way1Dirty_26 = _RAND_794[0:0];
  _RAND_795 = {1{`RANDOM}};
  way1Dirty_27 = _RAND_795[0:0];
  _RAND_796 = {1{`RANDOM}};
  way1Dirty_28 = _RAND_796[0:0];
  _RAND_797 = {1{`RANDOM}};
  way1Dirty_29 = _RAND_797[0:0];
  _RAND_798 = {1{`RANDOM}};
  way1Dirty_30 = _RAND_798[0:0];
  _RAND_799 = {1{`RANDOM}};
  way1Dirty_31 = _RAND_799[0:0];
  _RAND_800 = {1{`RANDOM}};
  way1Dirty_32 = _RAND_800[0:0];
  _RAND_801 = {1{`RANDOM}};
  way1Dirty_33 = _RAND_801[0:0];
  _RAND_802 = {1{`RANDOM}};
  way1Dirty_34 = _RAND_802[0:0];
  _RAND_803 = {1{`RANDOM}};
  way1Dirty_35 = _RAND_803[0:0];
  _RAND_804 = {1{`RANDOM}};
  way1Dirty_36 = _RAND_804[0:0];
  _RAND_805 = {1{`RANDOM}};
  way1Dirty_37 = _RAND_805[0:0];
  _RAND_806 = {1{`RANDOM}};
  way1Dirty_38 = _RAND_806[0:0];
  _RAND_807 = {1{`RANDOM}};
  way1Dirty_39 = _RAND_807[0:0];
  _RAND_808 = {1{`RANDOM}};
  way1Dirty_40 = _RAND_808[0:0];
  _RAND_809 = {1{`RANDOM}};
  way1Dirty_41 = _RAND_809[0:0];
  _RAND_810 = {1{`RANDOM}};
  way1Dirty_42 = _RAND_810[0:0];
  _RAND_811 = {1{`RANDOM}};
  way1Dirty_43 = _RAND_811[0:0];
  _RAND_812 = {1{`RANDOM}};
  way1Dirty_44 = _RAND_812[0:0];
  _RAND_813 = {1{`RANDOM}};
  way1Dirty_45 = _RAND_813[0:0];
  _RAND_814 = {1{`RANDOM}};
  way1Dirty_46 = _RAND_814[0:0];
  _RAND_815 = {1{`RANDOM}};
  way1Dirty_47 = _RAND_815[0:0];
  _RAND_816 = {1{`RANDOM}};
  way1Dirty_48 = _RAND_816[0:0];
  _RAND_817 = {1{`RANDOM}};
  way1Dirty_49 = _RAND_817[0:0];
  _RAND_818 = {1{`RANDOM}};
  way1Dirty_50 = _RAND_818[0:0];
  _RAND_819 = {1{`RANDOM}};
  way1Dirty_51 = _RAND_819[0:0];
  _RAND_820 = {1{`RANDOM}};
  way1Dirty_52 = _RAND_820[0:0];
  _RAND_821 = {1{`RANDOM}};
  way1Dirty_53 = _RAND_821[0:0];
  _RAND_822 = {1{`RANDOM}};
  way1Dirty_54 = _RAND_822[0:0];
  _RAND_823 = {1{`RANDOM}};
  way1Dirty_55 = _RAND_823[0:0];
  _RAND_824 = {1{`RANDOM}};
  way1Dirty_56 = _RAND_824[0:0];
  _RAND_825 = {1{`RANDOM}};
  way1Dirty_57 = _RAND_825[0:0];
  _RAND_826 = {1{`RANDOM}};
  way1Dirty_58 = _RAND_826[0:0];
  _RAND_827 = {1{`RANDOM}};
  way1Dirty_59 = _RAND_827[0:0];
  _RAND_828 = {1{`RANDOM}};
  way1Dirty_60 = _RAND_828[0:0];
  _RAND_829 = {1{`RANDOM}};
  way1Dirty_61 = _RAND_829[0:0];
  _RAND_830 = {1{`RANDOM}};
  way1Dirty_62 = _RAND_830[0:0];
  _RAND_831 = {1{`RANDOM}};
  way1Dirty_63 = _RAND_831[0:0];
  _RAND_832 = {1{`RANDOM}};
  way1Dirty_64 = _RAND_832[0:0];
  _RAND_833 = {1{`RANDOM}};
  way1Dirty_65 = _RAND_833[0:0];
  _RAND_834 = {1{`RANDOM}};
  way1Dirty_66 = _RAND_834[0:0];
  _RAND_835 = {1{`RANDOM}};
  way1Dirty_67 = _RAND_835[0:0];
  _RAND_836 = {1{`RANDOM}};
  way1Dirty_68 = _RAND_836[0:0];
  _RAND_837 = {1{`RANDOM}};
  way1Dirty_69 = _RAND_837[0:0];
  _RAND_838 = {1{`RANDOM}};
  way1Dirty_70 = _RAND_838[0:0];
  _RAND_839 = {1{`RANDOM}};
  way1Dirty_71 = _RAND_839[0:0];
  _RAND_840 = {1{`RANDOM}};
  way1Dirty_72 = _RAND_840[0:0];
  _RAND_841 = {1{`RANDOM}};
  way1Dirty_73 = _RAND_841[0:0];
  _RAND_842 = {1{`RANDOM}};
  way1Dirty_74 = _RAND_842[0:0];
  _RAND_843 = {1{`RANDOM}};
  way1Dirty_75 = _RAND_843[0:0];
  _RAND_844 = {1{`RANDOM}};
  way1Dirty_76 = _RAND_844[0:0];
  _RAND_845 = {1{`RANDOM}};
  way1Dirty_77 = _RAND_845[0:0];
  _RAND_846 = {1{`RANDOM}};
  way1Dirty_78 = _RAND_846[0:0];
  _RAND_847 = {1{`RANDOM}};
  way1Dirty_79 = _RAND_847[0:0];
  _RAND_848 = {1{`RANDOM}};
  way1Dirty_80 = _RAND_848[0:0];
  _RAND_849 = {1{`RANDOM}};
  way1Dirty_81 = _RAND_849[0:0];
  _RAND_850 = {1{`RANDOM}};
  way1Dirty_82 = _RAND_850[0:0];
  _RAND_851 = {1{`RANDOM}};
  way1Dirty_83 = _RAND_851[0:0];
  _RAND_852 = {1{`RANDOM}};
  way1Dirty_84 = _RAND_852[0:0];
  _RAND_853 = {1{`RANDOM}};
  way1Dirty_85 = _RAND_853[0:0];
  _RAND_854 = {1{`RANDOM}};
  way1Dirty_86 = _RAND_854[0:0];
  _RAND_855 = {1{`RANDOM}};
  way1Dirty_87 = _RAND_855[0:0];
  _RAND_856 = {1{`RANDOM}};
  way1Dirty_88 = _RAND_856[0:0];
  _RAND_857 = {1{`RANDOM}};
  way1Dirty_89 = _RAND_857[0:0];
  _RAND_858 = {1{`RANDOM}};
  way1Dirty_90 = _RAND_858[0:0];
  _RAND_859 = {1{`RANDOM}};
  way1Dirty_91 = _RAND_859[0:0];
  _RAND_860 = {1{`RANDOM}};
  way1Dirty_92 = _RAND_860[0:0];
  _RAND_861 = {1{`RANDOM}};
  way1Dirty_93 = _RAND_861[0:0];
  _RAND_862 = {1{`RANDOM}};
  way1Dirty_94 = _RAND_862[0:0];
  _RAND_863 = {1{`RANDOM}};
  way1Dirty_95 = _RAND_863[0:0];
  _RAND_864 = {1{`RANDOM}};
  way1Dirty_96 = _RAND_864[0:0];
  _RAND_865 = {1{`RANDOM}};
  way1Dirty_97 = _RAND_865[0:0];
  _RAND_866 = {1{`RANDOM}};
  way1Dirty_98 = _RAND_866[0:0];
  _RAND_867 = {1{`RANDOM}};
  way1Dirty_99 = _RAND_867[0:0];
  _RAND_868 = {1{`RANDOM}};
  way1Dirty_100 = _RAND_868[0:0];
  _RAND_869 = {1{`RANDOM}};
  way1Dirty_101 = _RAND_869[0:0];
  _RAND_870 = {1{`RANDOM}};
  way1Dirty_102 = _RAND_870[0:0];
  _RAND_871 = {1{`RANDOM}};
  way1Dirty_103 = _RAND_871[0:0];
  _RAND_872 = {1{`RANDOM}};
  way1Dirty_104 = _RAND_872[0:0];
  _RAND_873 = {1{`RANDOM}};
  way1Dirty_105 = _RAND_873[0:0];
  _RAND_874 = {1{`RANDOM}};
  way1Dirty_106 = _RAND_874[0:0];
  _RAND_875 = {1{`RANDOM}};
  way1Dirty_107 = _RAND_875[0:0];
  _RAND_876 = {1{`RANDOM}};
  way1Dirty_108 = _RAND_876[0:0];
  _RAND_877 = {1{`RANDOM}};
  way1Dirty_109 = _RAND_877[0:0];
  _RAND_878 = {1{`RANDOM}};
  way1Dirty_110 = _RAND_878[0:0];
  _RAND_879 = {1{`RANDOM}};
  way1Dirty_111 = _RAND_879[0:0];
  _RAND_880 = {1{`RANDOM}};
  way1Dirty_112 = _RAND_880[0:0];
  _RAND_881 = {1{`RANDOM}};
  way1Dirty_113 = _RAND_881[0:0];
  _RAND_882 = {1{`RANDOM}};
  way1Dirty_114 = _RAND_882[0:0];
  _RAND_883 = {1{`RANDOM}};
  way1Dirty_115 = _RAND_883[0:0];
  _RAND_884 = {1{`RANDOM}};
  way1Dirty_116 = _RAND_884[0:0];
  _RAND_885 = {1{`RANDOM}};
  way1Dirty_117 = _RAND_885[0:0];
  _RAND_886 = {1{`RANDOM}};
  way1Dirty_118 = _RAND_886[0:0];
  _RAND_887 = {1{`RANDOM}};
  way1Dirty_119 = _RAND_887[0:0];
  _RAND_888 = {1{`RANDOM}};
  way1Dirty_120 = _RAND_888[0:0];
  _RAND_889 = {1{`RANDOM}};
  way1Dirty_121 = _RAND_889[0:0];
  _RAND_890 = {1{`RANDOM}};
  way1Dirty_122 = _RAND_890[0:0];
  _RAND_891 = {1{`RANDOM}};
  way1Dirty_123 = _RAND_891[0:0];
  _RAND_892 = {1{`RANDOM}};
  way1Dirty_124 = _RAND_892[0:0];
  _RAND_893 = {1{`RANDOM}};
  way1Dirty_125 = _RAND_893[0:0];
  _RAND_894 = {1{`RANDOM}};
  way1Dirty_126 = _RAND_894[0:0];
  _RAND_895 = {1{`RANDOM}};
  way1Dirty_127 = _RAND_895[0:0];
  _RAND_896 = {1{`RANDOM}};
  state = _RAND_896[2:0];
  _RAND_897 = {1{`RANDOM}};
  cacheWriteEn_REG = _RAND_897[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AxiLite2Axi(
  input          clock,
  input          reset,
  input          io_out_aw_ready,
  output         io_out_aw_valid,
  output [31:0]  io_out_aw_bits_addr,
  input          io_out_w_ready,
  output         io_out_w_valid,
  output [63:0]  io_out_w_bits_data,
  output [7:0]   io_out_w_bits_strb,
  output         io_out_w_bits_last,
  output         io_out_b_ready,
  input          io_out_b_valid,
  input          io_out_ar_ready,
  output         io_out_ar_valid,
  output [31:0]  io_out_ar_bits_addr,
  output         io_out_r_ready,
  input          io_out_r_valid,
  input  [63:0]  io_out_r_bits_data,
  input          io_out_r_bits_last,
  input          io_imem_inst_valid,
  output         io_imem_inst_ready,
  input  [31:0]  io_imem_inst_addr,
  output [127:0] io_imem_inst_read,
  input          io_dmem_data_valid,
  output         io_dmem_data_ready,
  input          io_dmem_data_req,
  input  [31:0]  io_dmem_data_addr,
  input  [7:0]   io_dmem_data_strb,
  output [127:0] io_dmem_data_read,
  input  [127:0] io_dmem_data_write
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  wire  data_ren = io_dmem_data_valid & ~io_dmem_data_req; // @[Axi.scala 29:30]
  wire  data_wen = io_dmem_data_valid & io_dmem_data_req; // @[Axi.scala 30:30]
  wire  ar_hs = io_out_ar_ready & io_out_ar_valid; // @[Axi.scala 32:28]
  wire  r_hs = io_out_r_valid & io_out_r_ready; // @[Axi.scala 33:26]
  wire  aw_hs = io_out_aw_ready & io_out_aw_valid; // @[Axi.scala 34:28]
  wire  w_hs = io_out_w_ready & io_out_w_valid; // @[Axi.scala 35:26]
  wire  b_hs = io_out_b_valid & io_out_b_ready; // @[Axi.scala 36:26]
  wire  r_done = r_hs & io_out_r_bits_last; // @[Axi.scala 38:21]
  wire  w_done = b_hs & io_out_w_bits_last; // @[Axi.scala 39:21]
  reg [2:0] r_state; // @[Axi.scala 43:24]
  reg [2:0] w_state; // @[Axi.scala 44:24]
  wire [2:0] _GEN_3 = r_done ? 3'h3 : r_state; // @[Axi.scala 63:20 64:17 43:24]
  wire [2:0] _GEN_4 = data_ren ? 3'h4 : 3'h0; // @[Axi.scala 68:23 69:17 72:17]
  wire [2:0] _GEN_5 = ar_hs ? 3'h5 : r_state; // @[Axi.scala 77:20 78:17 43:24]
  wire [2:0] _GEN_6 = r_done ? 3'h6 : r_state; // @[Axi.scala 82:21 83:17 43:24]
  wire [2:0] _GEN_7 = 3'h6 == r_state ? 3'h0 : r_state; // @[Axi.scala 49:20 87:15 43:24]
  wire [2:0] _GEN_8 = 3'h5 == r_state ? _GEN_6 : _GEN_7; // @[Axi.scala 49:20]
  wire [2:0] _GEN_9 = 3'h4 == r_state ? _GEN_5 : _GEN_8; // @[Axi.scala 49:20]
  wire [2:0] _GEN_10 = 3'h3 == r_state ? _GEN_4 : _GEN_9; // @[Axi.scala 49:20]
  wire [2:0] _GEN_16 = w_hs ? 3'h3 : w_state; // @[Axi.scala 105:18 106:17 44:24]
  wire [2:0] _GEN_17 = w_done ? 3'h4 : w_state; // @[Axi.scala 110:20 111:17 44:24]
  wire [2:0] _GEN_18 = 3'h4 == w_state ? 3'h0 : w_state; // @[Axi.scala 115:15 93:20 44:24]
  wire [2:0] _GEN_19 = 3'h3 == w_state ? _GEN_17 : _GEN_18; // @[Axi.scala 93:20]
  reg  data_ok; // @[Axi.scala 119:24]
  wire  _T_12 = w_state == 3'h4; // @[Axi.scala 120:29]
  wire  _GEN_23 = ~data_wen ? 1'h0 : data_ok; // @[Axi.scala 123:25 124:13 119:24]
  wire  _GEN_24 = data_wen & w_state == 3'h4 | _GEN_23; // @[Axi.scala 120:46 121:13]
  wire  _axi_addr_T = r_state == 3'h1; // @[Axi.scala 127:30]
  wire [31:0] _axi_addr_T_1 = io_imem_inst_addr & 32'hfffffff0; // @[Axi.scala 127:63]
  wire  _axi_addr_T_2 = r_state == 3'h4; // @[Axi.scala 128:31]
  wire [31:0] _axi_addr_T_3 = io_dmem_data_addr & 32'hfffffff0; // @[Axi.scala 128:64]
  wire [31:0] _axi_addr_T_4 = r_state == 3'h4 ? _axi_addr_T_3 : 32'h0; // @[Axi.scala 128:22]
  wire [31:0] _axi_waddr_T_1 = {io_dmem_data_addr[31:4],4'h8}; // @[Cat.scala 31:58]
  wire [31:0] _GEN_33 = io_dmem_data_addr % 32'h10; // @[Axi.scala 150:38]
  wire  lowDateEn = _GEN_33[4:0] < 5'h8; // @[Axi.scala 150:46]
  wire [7:0] strb_h = ~lowDateEn ? io_dmem_data_strb : 8'h0; // @[Axi.scala 151:19]
  wire [7:0] strb_l = lowDateEn ? io_dmem_data_strb : 8'h0; // @[Axi.scala 152:19]
  reg [63:0] inst_read_h; // @[Axi.scala 178:28]
  reg [63:0] inst_read_l; // @[Axi.scala 179:28]
  reg [63:0] data_read_h; // @[Axi.scala 180:28]
  reg [63:0] data_read_l; // @[Axi.scala 181:28]
  wire [127:0] dmemData = {data_read_h,data_read_l}; // @[Cat.scala 31:58]
  wire [8:0] _io_dmem_data_read_T = _GEN_33[4:0] * 4'h8; // @[Axi.scala 197:42]
  assign io_out_aw_valid = w_state == 3'h1; // @[Axi.scala 154:34]
  assign io_out_aw_bits_addr = data_ok ? _axi_waddr_T_1 : _axi_addr_T_3; // @[Axi.scala 149:22]
  assign io_out_w_valid = w_state == 3'h2; // @[Axi.scala 167:34]
  assign io_out_w_bits_data = data_ok ? io_dmem_data_write[127:64] : io_dmem_data_write[63:0]; // @[Axi.scala 168:29]
  assign io_out_w_bits_strb = data_ok ? strb_h : strb_l; // @[Axi.scala 169:29]
  assign io_out_w_bits_last = 1'h1; // @[Axi.scala 170:23]
  assign io_out_b_ready = 1'h1; // @[Axi.scala 172:23]
  assign io_out_ar_valid = _axi_addr_T | _axi_addr_T_2; // @[Axi.scala 130:44]
  assign io_out_ar_bits_addr = r_state == 3'h1 ? _axi_addr_T_1 : _axi_addr_T_4; // @[Axi.scala 127:21]
  assign io_out_r_ready = 1'h1; // @[Axi.scala 143:15]
  assign io_imem_inst_ready = r_state == 3'h3; // @[Axi.scala 175:30]
  assign io_imem_inst_read = {inst_read_h,inst_read_l}; // @[Cat.scala 31:58]
  assign io_dmem_data_ready = r_state == 3'h6 | _T_12 & data_ok; // @[Axi.scala 176:47]
  assign io_dmem_data_read = dmemData >> _io_dmem_data_read_T; // @[Axi.scala 197:29]
  always @(posedge clock) begin
    if (reset) begin // @[Axi.scala 43:24]
      r_state <= 3'h0; // @[Axi.scala 43:24]
    end else if (3'h0 == r_state) begin // @[Axi.scala 49:20]
      if (io_imem_inst_valid) begin // @[Axi.scala 51:22]
        r_state <= 3'h1; // @[Axi.scala 52:17]
      end else if (data_ren) begin // @[Axi.scala 53:30]
        r_state <= 3'h4; // @[Axi.scala 54:17]
      end
    end else if (3'h1 == r_state) begin // @[Axi.scala 49:20]
      if (ar_hs) begin // @[Axi.scala 58:19]
        r_state <= 3'h2; // @[Axi.scala 59:17]
      end
    end else if (3'h2 == r_state) begin // @[Axi.scala 49:20]
      r_state <= _GEN_3;
    end else begin
      r_state <= _GEN_10;
    end
    if (reset) begin // @[Axi.scala 44:24]
      w_state <= 3'h0; // @[Axi.scala 44:24]
    end else if (3'h0 == w_state) begin // @[Axi.scala 93:20]
      if (data_wen) begin // @[Axi.scala 95:22]
        w_state <= 3'h1; // @[Axi.scala 96:17]
      end
    end else if (3'h1 == w_state) begin // @[Axi.scala 93:20]
      if (aw_hs) begin // @[Axi.scala 100:19]
        w_state <= 3'h2; // @[Axi.scala 101:17]
      end
    end else if (3'h2 == w_state) begin // @[Axi.scala 93:20]
      w_state <= _GEN_16;
    end else begin
      w_state <= _GEN_19;
    end
    if (reset) begin // @[Axi.scala 119:24]
      data_ok <= 1'h0; // @[Axi.scala 119:24]
    end else begin
      data_ok <= _GEN_24;
    end
    if (reset) begin // @[Axi.scala 178:28]
      inst_read_h <= 64'h0; // @[Axi.scala 178:28]
    end else if (r_hs) begin // @[Axi.scala 183:15]
      if (io_out_r_bits_last) begin // @[Axi.scala 184:28]
        inst_read_h <= io_out_r_bits_data; // @[Axi.scala 185:19]
      end
    end
    if (reset) begin // @[Axi.scala 179:28]
      inst_read_l <= 64'h0; // @[Axi.scala 179:28]
    end else if (r_hs) begin // @[Axi.scala 183:15]
      if (!(io_out_r_bits_last)) begin // @[Axi.scala 184:28]
        inst_read_l <= io_out_r_bits_data; // @[Axi.scala 189:19]
      end
    end
    if (reset) begin // @[Axi.scala 180:28]
      data_read_h <= 64'h0; // @[Axi.scala 180:28]
    end else if (r_hs) begin // @[Axi.scala 183:15]
      if (io_out_r_bits_last) begin // @[Axi.scala 184:28]
        data_read_h <= io_out_r_bits_data; // @[Axi.scala 186:19]
      end
    end
    if (reset) begin // @[Axi.scala 181:28]
      data_read_l <= 64'h0; // @[Axi.scala 181:28]
    end else if (r_hs) begin // @[Axi.scala 183:15]
      if (!(io_out_r_bits_last)) begin // @[Axi.scala 184:28]
        data_read_l <= io_out_r_bits_data; // @[Axi.scala 190:19]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r_state = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  w_state = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  data_ok = _RAND_2[0:0];
  _RAND_3 = {2{`RANDOM}};
  inst_read_h = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  inst_read_l = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  data_read_h = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  data_read_l = _RAND_6[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SimTop(
  input         clock,
  input         reset,
  input  [63:0] io_logCtrl_log_begin,
  input  [63:0] io_logCtrl_log_end,
  input  [63:0] io_logCtrl_log_level,
  input         io_perfInfo_clean,
  input         io_perfInfo_dump,
  output        io_uart_out_valid,
  output [7:0]  io_uart_out_ch,
  output        io_uart_in_valid,
  input  [7:0]  io_uart_in_ch,
  input         io_memAXI_0_aw_ready,
  output        io_memAXI_0_aw_valid,
  output [31:0] io_memAXI_0_aw_bits_addr,
  output [2:0]  io_memAXI_0_aw_bits_prot,
  output [3:0]  io_memAXI_0_aw_bits_id,
  output        io_memAXI_0_aw_bits_user,
  output [7:0]  io_memAXI_0_aw_bits_len,
  output [2:0]  io_memAXI_0_aw_bits_size,
  output [1:0]  io_memAXI_0_aw_bits_burst,
  output        io_memAXI_0_aw_bits_lock,
  output [3:0]  io_memAXI_0_aw_bits_cache,
  output [3:0]  io_memAXI_0_aw_bits_qos,
  input         io_memAXI_0_w_ready,
  output        io_memAXI_0_w_valid,
  output [63:0] io_memAXI_0_w_bits_data[3:0],
  output [7:0]  io_memAXI_0_w_bits_strb,
  output        io_memAXI_0_w_bits_last,
  output        io_memAXI_0_b_ready,
  input         io_memAXI_0_b_valid,
  input  [1:0]  io_memAXI_0_b_bits_resp,
  input  [3:0]  io_memAXI_0_b_bits_id,
  input         io_memAXI_0_b_bits_user,
  input         io_memAXI_0_ar_ready,
  output        io_memAXI_0_ar_valid,
  output [31:0] io_memAXI_0_ar_bits_addr,
  output [2:0]  io_memAXI_0_ar_bits_prot,
  output [3:0]  io_memAXI_0_ar_bits_id,
  output        io_memAXI_0_ar_bits_user,
  output [7:0]  io_memAXI_0_ar_bits_len,
  output [2:0]  io_memAXI_0_ar_bits_size,
  output [1:0]  io_memAXI_0_ar_bits_burst,
  output        io_memAXI_0_ar_bits_lock,
  output [3:0]  io_memAXI_0_ar_bits_cache,
  output [3:0]  io_memAXI_0_ar_bits_qos,
  output        io_memAXI_0_r_ready,
  input         io_memAXI_0_r_valid,
  input  [1:0]  io_memAXI_0_r_bits_resp,
  input  [63:0] io_memAXI_0_r_bits_data[3:0],
  input  [3:0]  io_memAXI_0_r_bits_id,
  input         io_memAXI_0_r_bits_user,
  input         io_memAXI_0_r_bits_last
);
  wire  core_clock; // @[SimTop.scala 18:20]
  wire  core_reset; // @[SimTop.scala 18:20]
  wire  core_io_imem_inst_valid; // @[SimTop.scala 18:20]
  wire  core_io_imem_inst_ready; // @[SimTop.scala 18:20]
  wire [31:0] core_io_imem_inst_addr; // @[SimTop.scala 18:20]
  wire [31:0] core_io_imem_inst_read; // @[SimTop.scala 18:20]
  wire  core_io_dmem_data_valid; // @[SimTop.scala 18:20]
  wire  core_io_dmem_data_ready; // @[SimTop.scala 18:20]
  wire  core_io_dmem_data_req; // @[SimTop.scala 18:20]
  wire [31:0] core_io_dmem_data_addr; // @[SimTop.scala 18:20]
  wire [1:0] core_io_dmem_data_size; // @[SimTop.scala 18:20]
  wire [7:0] core_io_dmem_data_strb; // @[SimTop.scala 18:20]
  wire [63:0] core_io_dmem_data_read; // @[SimTop.scala 18:20]
  wire [127:0] core_io_dmem_data_write; // @[SimTop.scala 18:20]
  wire  icache_clock; // @[SimTop.scala 19:22]
  wire  icache_reset; // @[SimTop.scala 19:22]
  wire  icache_io_imem_inst_valid; // @[SimTop.scala 19:22]
  wire  icache_io_imem_inst_ready; // @[SimTop.scala 19:22]
  wire [31:0] icache_io_imem_inst_addr; // @[SimTop.scala 19:22]
  wire [31:0] icache_io_imem_inst_read; // @[SimTop.scala 19:22]
  wire  icache_io_out_inst_valid; // @[SimTop.scala 19:22]
  wire  icache_io_out_inst_ready; // @[SimTop.scala 19:22]
  wire [31:0] icache_io_out_inst_addr; // @[SimTop.scala 19:22]
  wire [127:0] icache_io_out_inst_read; // @[SimTop.scala 19:22]
  wire  dcache_clock; // @[SimTop.scala 20:22]
  wire  dcache_reset; // @[SimTop.scala 20:22]
  wire  dcache_io_dmem_data_valid; // @[SimTop.scala 20:22]
  wire  dcache_io_dmem_data_ready; // @[SimTop.scala 20:22]
  wire  dcache_io_dmem_data_req; // @[SimTop.scala 20:22]
  wire [31:0] dcache_io_dmem_data_addr; // @[SimTop.scala 20:22]
  wire [1:0] dcache_io_dmem_data_size; // @[SimTop.scala 20:22]
  wire [7:0] dcache_io_dmem_data_strb; // @[SimTop.scala 20:22]
  wire [63:0] dcache_io_dmem_data_read; // @[SimTop.scala 20:22]
  wire [127:0] dcache_io_dmem_data_write; // @[SimTop.scala 20:22]
  wire  dcache_io_out_data_valid; // @[SimTop.scala 20:22]
  wire  dcache_io_out_data_ready; // @[SimTop.scala 20:22]
  wire  dcache_io_out_data_req; // @[SimTop.scala 20:22]
  wire [31:0] dcache_io_out_data_addr; // @[SimTop.scala 20:22]
  wire [7:0] dcache_io_out_data_strb; // @[SimTop.scala 20:22]
  wire [127:0] dcache_io_out_data_read; // @[SimTop.scala 20:22]
  wire [127:0] dcache_io_out_data_write; // @[SimTop.scala 20:22]
  wire  top_clock; // @[SimTop.scala 23:19]
  wire  top_reset; // @[SimTop.scala 23:19]
  wire  top_io_out_aw_ready; // @[SimTop.scala 23:19]
  wire  top_io_out_aw_valid; // @[SimTop.scala 23:19]
  wire [31:0] top_io_out_aw_bits_addr; // @[SimTop.scala 23:19]
  wire  top_io_out_w_ready; // @[SimTop.scala 23:19]
  wire  top_io_out_w_valid; // @[SimTop.scala 23:19]
  wire [63:0] top_io_out_w_bits_data; // @[SimTop.scala 23:19]
  wire [7:0] top_io_out_w_bits_strb; // @[SimTop.scala 23:19]
  wire  top_io_out_w_bits_last; // @[SimTop.scala 23:19]
  wire  top_io_out_b_ready; // @[SimTop.scala 23:19]
  wire  top_io_out_b_valid; // @[SimTop.scala 23:19]
  wire  top_io_out_ar_ready; // @[SimTop.scala 23:19]
  wire  top_io_out_ar_valid; // @[SimTop.scala 23:19]
  wire [31:0] top_io_out_ar_bits_addr; // @[SimTop.scala 23:19]
  wire  top_io_out_r_ready; // @[SimTop.scala 23:19]
  wire  top_io_out_r_valid; // @[SimTop.scala 23:19]
  wire [63:0] top_io_out_r_bits_data; // @[SimTop.scala 23:19]
  wire  top_io_out_r_bits_last; // @[SimTop.scala 23:19]
  wire  top_io_imem_inst_valid; // @[SimTop.scala 23:19]
  wire  top_io_imem_inst_ready; // @[SimTop.scala 23:19]
  wire [31:0] top_io_imem_inst_addr; // @[SimTop.scala 23:19]
  wire [127:0] top_io_imem_inst_read; // @[SimTop.scala 23:19]
  wire  top_io_dmem_data_valid; // @[SimTop.scala 23:19]
  wire  top_io_dmem_data_ready; // @[SimTop.scala 23:19]
  wire  top_io_dmem_data_req; // @[SimTop.scala 23:19]
  wire [31:0] top_io_dmem_data_addr; // @[SimTop.scala 23:19]
  wire [7:0] top_io_dmem_data_strb; // @[SimTop.scala 23:19]
  wire [127:0] top_io_dmem_data_read; // @[SimTop.scala 23:19]
  wire [127:0] top_io_dmem_data_write; // @[SimTop.scala 23:19]
  Core core ( // @[SimTop.scala 18:20]
    .clock(core_clock),
    .reset(core_reset),
    .io_imem_inst_valid(core_io_imem_inst_valid),
    .io_imem_inst_ready(core_io_imem_inst_ready),
    .io_imem_inst_addr(core_io_imem_inst_addr),
    .io_imem_inst_read(core_io_imem_inst_read),
    .io_dmem_data_valid(core_io_dmem_data_valid),
    .io_dmem_data_ready(core_io_dmem_data_ready),
    .io_dmem_data_req(core_io_dmem_data_req),
    .io_dmem_data_addr(core_io_dmem_data_addr),
    .io_dmem_data_size(core_io_dmem_data_size),
    .io_dmem_data_strb(core_io_dmem_data_strb),
    .io_dmem_data_read(core_io_dmem_data_read),
    .io_dmem_data_write(core_io_dmem_data_write)
  );
  ICache icache ( // @[SimTop.scala 19:22]
    .clock(icache_clock),
    .reset(icache_reset),
    .io_imem_inst_valid(icache_io_imem_inst_valid),
    .io_imem_inst_ready(icache_io_imem_inst_ready),
    .io_imem_inst_addr(icache_io_imem_inst_addr),
    .io_imem_inst_read(icache_io_imem_inst_read),
    .io_out_inst_valid(icache_io_out_inst_valid),
    .io_out_inst_ready(icache_io_out_inst_ready),
    .io_out_inst_addr(icache_io_out_inst_addr),
    .io_out_inst_read(icache_io_out_inst_read)
  );
  DCache dcache ( // @[SimTop.scala 20:22]
    .clock(dcache_clock),
    .reset(dcache_reset),
    .io_dmem_data_valid(dcache_io_dmem_data_valid),
    .io_dmem_data_ready(dcache_io_dmem_data_ready),
    .io_dmem_data_req(dcache_io_dmem_data_req),
    .io_dmem_data_addr(dcache_io_dmem_data_addr),
    .io_dmem_data_size(dcache_io_dmem_data_size),
    .io_dmem_data_strb(dcache_io_dmem_data_strb),
    .io_dmem_data_read(dcache_io_dmem_data_read),
    .io_dmem_data_write(dcache_io_dmem_data_write),
    .io_out_data_valid(dcache_io_out_data_valid),
    .io_out_data_ready(dcache_io_out_data_ready),
    .io_out_data_req(dcache_io_out_data_req),
    .io_out_data_addr(dcache_io_out_data_addr),
    .io_out_data_strb(dcache_io_out_data_strb),
    .io_out_data_read(dcache_io_out_data_read),
    .io_out_data_write(dcache_io_out_data_write)
  );
  AxiLite2Axi top ( // @[SimTop.scala 23:19]
    .clock(top_clock),
    .reset(top_reset),
    .io_out_aw_ready(top_io_out_aw_ready),
    .io_out_aw_valid(top_io_out_aw_valid),
    .io_out_aw_bits_addr(top_io_out_aw_bits_addr),
    .io_out_w_ready(top_io_out_w_ready),
    .io_out_w_valid(top_io_out_w_valid),
    .io_out_w_bits_data(top_io_out_w_bits_data),
    .io_out_w_bits_strb(top_io_out_w_bits_strb),
    .io_out_w_bits_last(top_io_out_w_bits_last),
    .io_out_b_ready(top_io_out_b_ready),
    .io_out_b_valid(top_io_out_b_valid),
    .io_out_ar_ready(top_io_out_ar_ready),
    .io_out_ar_valid(top_io_out_ar_valid),
    .io_out_ar_bits_addr(top_io_out_ar_bits_addr),
    .io_out_r_ready(top_io_out_r_ready),
    .io_out_r_valid(top_io_out_r_valid),
    .io_out_r_bits_data(top_io_out_r_bits_data),
    .io_out_r_bits_last(top_io_out_r_bits_last),
    .io_imem_inst_valid(top_io_imem_inst_valid),
    .io_imem_inst_ready(top_io_imem_inst_ready),
    .io_imem_inst_addr(top_io_imem_inst_addr),
    .io_imem_inst_read(top_io_imem_inst_read),
    .io_dmem_data_valid(top_io_dmem_data_valid),
    .io_dmem_data_ready(top_io_dmem_data_ready),
    .io_dmem_data_req(top_io_dmem_data_req),
    .io_dmem_data_addr(top_io_dmem_data_addr),
    .io_dmem_data_strb(top_io_dmem_data_strb),
    .io_dmem_data_read(top_io_dmem_data_read),
    .io_dmem_data_write(top_io_dmem_data_write)
  );
  assign io_uart_out_valid = 1'h0; // @[SimTop.scala 41:21]
  assign io_uart_out_ch = 8'h0; // @[SimTop.scala 42:18]
  assign io_uart_in_valid = 1'h0; // @[SimTop.scala 43:20]
  assign io_memAXI_0_aw_valid = top_io_out_aw_valid; // @[SimTop.scala 32:18]
  assign io_memAXI_0_aw_bits_addr = top_io_out_aw_bits_addr; // @[SimTop.scala 32:18]
  assign io_memAXI_0_aw_bits_prot = 3'h0; // @[SimTop.scala 32:18]
  assign io_memAXI_0_aw_bits_id = 4'h0; // @[SimTop.scala 32:18]
  assign io_memAXI_0_aw_bits_user = 1'h0; // @[SimTop.scala 32:18]
  assign io_memAXI_0_aw_bits_len = 8'h0; // @[SimTop.scala 32:18]
  assign io_memAXI_0_aw_bits_size = 3'h3; // @[SimTop.scala 32:18]
  assign io_memAXI_0_aw_bits_burst = 2'h1; // @[SimTop.scala 32:18]
  assign io_memAXI_0_aw_bits_lock = 1'h0; // @[SimTop.scala 32:18]
  assign io_memAXI_0_aw_bits_cache = 4'h2; // @[SimTop.scala 32:18]
  assign io_memAXI_0_aw_bits_qos = 4'h0; // @[SimTop.scala 32:18]
  assign io_memAXI_0_w_valid = top_io_out_w_valid; // @[SimTop.scala 33:18]
  assign io_memAXI_0_w_bits_data[0] = top_io_out_w_bits_data; // @[SimTop.scala 33:18]
  assign io_memAXI_0_w_bits_strb = top_io_out_w_bits_strb; // @[SimTop.scala 33:18]
  assign io_memAXI_0_w_bits_last = 1'h1; // @[SimTop.scala 33:18]
  assign io_memAXI_0_b_ready = 1'h1; // @[SimTop.scala 34:18]
  assign io_memAXI_0_ar_valid = top_io_out_ar_valid; // @[SimTop.scala 35:18]
  assign io_memAXI_0_ar_bits_addr = top_io_out_ar_bits_addr; // @[SimTop.scala 35:18]
  assign io_memAXI_0_ar_bits_prot = 3'h0; // @[SimTop.scala 35:18]
  assign io_memAXI_0_ar_bits_id = 4'h0; // @[SimTop.scala 35:18]
  assign io_memAXI_0_ar_bits_user = 1'h0; // @[SimTop.scala 35:18]
  assign io_memAXI_0_ar_bits_len = 8'h1; // @[SimTop.scala 35:18]
  assign io_memAXI_0_ar_bits_size = 3'h3; // @[SimTop.scala 35:18]
  assign io_memAXI_0_ar_bits_burst = 2'h1; // @[SimTop.scala 35:18]
  assign io_memAXI_0_ar_bits_lock = 1'h0; // @[SimTop.scala 35:18]
  assign io_memAXI_0_ar_bits_cache = 4'h2; // @[SimTop.scala 35:18]
  assign io_memAXI_0_ar_bits_qos = 4'h0; // @[SimTop.scala 35:18]
  assign io_memAXI_0_r_ready = 1'h1; // @[SimTop.scala 36:18]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_imem_inst_ready = icache_io_imem_inst_ready; // @[SimTop.scala 27:17]
  assign core_io_imem_inst_read = icache_io_imem_inst_read; // @[SimTop.scala 27:17]
  assign core_io_dmem_data_ready = dcache_io_dmem_data_ready; // @[SimTop.scala 29:17]
  assign core_io_dmem_data_read = dcache_io_dmem_data_read; // @[SimTop.scala 29:17]
  assign icache_clock = clock;
  assign icache_reset = reset;
  assign icache_io_imem_inst_valid = core_io_imem_inst_valid; // @[SimTop.scala 27:17]
  assign icache_io_imem_inst_addr = core_io_imem_inst_addr; // @[SimTop.scala 27:17]
  assign icache_io_out_inst_ready = top_io_imem_inst_ready; // @[SimTop.scala 28:17]
  assign icache_io_out_inst_read = top_io_imem_inst_read; // @[SimTop.scala 28:17]
  assign dcache_clock = clock;
  assign dcache_reset = reset;
  assign dcache_io_dmem_data_valid = core_io_dmem_data_valid; // @[SimTop.scala 29:17]
  assign dcache_io_dmem_data_req = core_io_dmem_data_req; // @[SimTop.scala 29:17]
  assign dcache_io_dmem_data_addr = core_io_dmem_data_addr; // @[SimTop.scala 29:17]
  assign dcache_io_dmem_data_size = core_io_dmem_data_size; // @[SimTop.scala 29:17]
  assign dcache_io_dmem_data_strb = core_io_dmem_data_strb; // @[SimTop.scala 29:17]
  assign dcache_io_dmem_data_write = core_io_dmem_data_write; // @[SimTop.scala 29:17]
  assign dcache_io_out_data_ready = top_io_dmem_data_ready; // @[SimTop.scala 30:17]
  assign dcache_io_out_data_read = top_io_dmem_data_read; // @[SimTop.scala 30:17]
  assign top_clock = clock;
  assign top_reset = reset;
  assign top_io_out_aw_ready = io_memAXI_0_aw_ready; // @[SimTop.scala 32:18]
  assign top_io_out_w_ready = io_memAXI_0_w_ready; // @[SimTop.scala 33:18]
  assign top_io_out_b_valid = io_memAXI_0_b_valid; // @[SimTop.scala 34:18]
  assign top_io_out_ar_ready = io_memAXI_0_ar_ready; // @[SimTop.scala 35:18]
  assign top_io_out_r_valid = io_memAXI_0_r_valid; // @[SimTop.scala 36:18]
  assign top_io_out_r_bits_data = io_memAXI_0_r_bits_data[0]; // @[SimTop.scala 36:18]
  assign top_io_out_r_bits_last = io_memAXI_0_r_bits_last; // @[SimTop.scala 36:18]
  assign top_io_imem_inst_valid = icache_io_out_inst_valid; // @[SimTop.scala 28:17]
  assign top_io_imem_inst_addr = icache_io_out_inst_addr; // @[SimTop.scala 28:17]
  assign top_io_dmem_data_valid = dcache_io_out_data_valid; // @[SimTop.scala 30:17]
  assign top_io_dmem_data_req = dcache_io_out_data_req; // @[SimTop.scala 30:17]
  assign top_io_dmem_data_addr = dcache_io_out_data_addr; // @[SimTop.scala 30:17]
  assign top_io_dmem_data_strb = dcache_io_out_data_strb; // @[SimTop.scala 30:17]
  assign top_io_dmem_data_write = dcache_io_out_data_write; // @[SimTop.scala 30:17]
endmodule
