module ImmGen(
  input  [31:0] io_inst,
  input  [2:0]  io_immOp,
  output [63:0] io_imm
);
  wire [51:0] _immType_0_T_2 = io_inst[31] ? 52'hfffffffffffff : 52'h0; // @[Bitwise.scala 74:12]
  wire [63:0] immType_0 = {_immType_0_T_2,io_inst[31:20]}; // @[ImmGen.scala 19:41]
  wire [31:0] _immType_1_T_2 = io_inst[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] immType_1 = {_immType_1_T_2,io_inst[31:12],12'h0}; // @[ImmGen.scala 20:59]
  wire [63:0] immType_2 = {_immType_0_T_2,io_inst[31:25],io_inst[11:7]}; // @[ImmGen.scala 21:59]
  wire [64:0] _immType_3_T_11 = {_immType_0_T_2,io_inst[31],io_inst[7],io_inst[30:25],io_inst[11:8],1'h0}; // @[ImmGen.scala 22:113]
  wire [42:0] _immType_4_T_2 = io_inst[31] ? 43'h7ffffffffff : 43'h0; // @[Bitwise.scala 74:12]
  wire [63:0] immType_4 = {_immType_4_T_2,io_inst[31],io_inst[19:12],io_inst[20],io_inst[30:21],1'h0}; // @[ImmGen.scala 23:113]
  wire [63:0] _GEN_1 = 3'h1 == io_immOp ? immType_1 : immType_0; // @[ImmGen.scala 25:{16,16}]
  wire [63:0] _GEN_2 = 3'h2 == io_immOp ? immType_2 : _GEN_1; // @[ImmGen.scala 25:{16,16}]
  wire [63:0] immType_3 = _immType_3_T_11[63:0]; // @[ImmGen.scala 17:21 22:16]
  wire [63:0] _GEN_3 = 3'h3 == io_immOp ? immType_3 : _GEN_2; // @[ImmGen.scala 25:{16,16}]
  wire [63:0] _GEN_4 = 3'h4 == io_immOp ? immType_4 : _GEN_3; // @[ImmGen.scala 25:{16,16}]
  assign io_imm = io_immOp > 3'h4 ? 64'h0 : _GEN_4; // @[ImmGen.scala 25:16]
endmodule
module minidec(
  input  [31:0] io_inst,
  output        io_rs1En,
  output [4:0]  io_rs1Addr,
  output        io_bjp,
  output        io_jal,
  output        io_jalr,
  output        io_bxx,
  output [63:0] io_imm
);
  wire [31:0] imm_io_inst; // @[minidec.scala 49:19]
  wire [2:0] imm_io_immOp; // @[minidec.scala 49:19]
  wire [63:0] imm_io_imm; // @[minidec.scala 49:19]
  wire [31:0] _jalr_T = io_inst & 32'h707f; // @[minidec.scala 26:19]
  wire  jalr = 32'h67 == _jalr_T; // @[minidec.scala 26:19]
  wire [31:0] _jal_T = io_inst & 32'h7f; // @[minidec.scala 27:18]
  wire  jal = 32'h6f == _jal_T; // @[minidec.scala 27:18]
  wire  jxx = jal | jalr; // @[minidec.scala 28:16]
  wire  beq = 32'h63 == _jalr_T; // @[minidec.scala 30:18]
  wire  bne = 32'h1063 == _jalr_T; // @[minidec.scala 31:18]
  wire  blt = 32'h4063 == _jalr_T; // @[minidec.scala 32:18]
  wire  bge = 32'h5063 == _jalr_T; // @[minidec.scala 33:18]
  wire  bltu = 32'h6063 == _jalr_T; // @[minidec.scala 34:19]
  wire  bgeu = 32'h7063 == _jalr_T; // @[minidec.scala 35:19]
  wire  bxx = beq | bne | blt | bge | bltu | bgeu; // @[minidec.scala 36:38]
  wire  rs1En = jalr | bxx; // @[minidec.scala 39:20]
  wire [2:0] _immOp_T = jalr ? 3'h0 : 3'h5; // @[minidec.scala 46:18]
  wire [2:0] _immOp_T_1 = bxx ? 3'h3 : _immOp_T; // @[minidec.scala 45:17]
  ImmGen imm ( // @[minidec.scala 49:19]
    .io_inst(imm_io_inst),
    .io_immOp(imm_io_immOp),
    .io_imm(imm_io_imm)
  );
  assign io_rs1En = jalr | bxx; // @[minidec.scala 39:20]
  assign io_rs1Addr = rs1En ? io_inst[19:15] : 5'h0; // @[minidec.scala 41:20]
  assign io_bjp = jxx | bxx; // @[minidec.scala 38:16]
  assign io_jal = 32'h6f == _jal_T; // @[minidec.scala 27:18]
  assign io_jalr = 32'h67 == _jalr_T; // @[minidec.scala 26:19]
  assign io_bxx = beq | bne | blt | bge | bltu | bgeu; // @[minidec.scala 36:38]
  assign io_imm = imm_io_imm; // @[minidec.scala 59:10]
  assign imm_io_inst = io_inst; // @[minidec.scala 50:15]
  assign imm_io_immOp = jal ? 3'h4 : _immOp_T_1; // @[minidec.scala 44:15]
endmodule
module bht(
  input         clock,
  input         reset,
  input         io_valid,
  input         io_fire,
  input  [31:0] io_pc,
  input         io_jal,
  input         io_jalr,
  input         io_bxx,
  input  [63:0] io_imm,
  input  [4:0]  io_rs1Addr,
  input  [63:0] io_rs1Data,
  input  [63:0] io_rs1x1Data,
  input         io_exeX1En,
  input  [63:0] io_exeAluRes,
  input         io_memX1En,
  input  [63:0] io_memAluRes,
  input         io_wbRdEn,
  input  [4:0]  io_wbRdAddr,
  input  [63:0] io_wbRdData,
  input         io_takenValid,
  input         io_takenValidJalr,
  input         io_takenMiss,
  input         io_exTakenPre,
  input  [31:0] io_takenPC,
  input  [31:0] io_nextPC,
  output        io_takenPre,
  output [31:0] io_takenPrePC,
  output        io_ready
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_645;
  reg [31:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_649;
  reg [31:0] _RAND_650;
  reg [31:0] _RAND_651;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
  reg [31:0] _RAND_654;
  reg [31:0] _RAND_655;
  reg [31:0] _RAND_656;
  reg [31:0] _RAND_657;
  reg [31:0] _RAND_658;
  reg [31:0] _RAND_659;
  reg [31:0] _RAND_660;
  reg [31:0] _RAND_661;
  reg [31:0] _RAND_662;
  reg [31:0] _RAND_663;
  reg [31:0] _RAND_664;
  reg [31:0] _RAND_665;
  reg [31:0] _RAND_666;
  reg [31:0] _RAND_667;
  reg [31:0] _RAND_668;
  reg [31:0] _RAND_669;
  reg [31:0] _RAND_670;
  reg [31:0] _RAND_671;
  reg [31:0] _RAND_672;
  reg [31:0] _RAND_673;
  reg [31:0] _RAND_674;
  reg [31:0] _RAND_675;
  reg [31:0] _RAND_676;
  reg [31:0] _RAND_677;
  reg [31:0] _RAND_678;
  reg [31:0] _RAND_679;
  reg [31:0] _RAND_680;
  reg [31:0] _RAND_681;
  reg [31:0] _RAND_682;
  reg [31:0] _RAND_683;
  reg [31:0] _RAND_684;
  reg [31:0] _RAND_685;
  reg [31:0] _RAND_686;
  reg [31:0] _RAND_687;
  reg [31:0] _RAND_688;
  reg [31:0] _RAND_689;
  reg [31:0] _RAND_690;
  reg [31:0] _RAND_691;
  reg [31:0] _RAND_692;
  reg [31:0] _RAND_693;
  reg [31:0] _RAND_694;
  reg [31:0] _RAND_695;
  reg [31:0] _RAND_696;
  reg [31:0] _RAND_697;
  reg [31:0] _RAND_698;
  reg [31:0] _RAND_699;
  reg [31:0] _RAND_700;
  reg [31:0] _RAND_701;
  reg [31:0] _RAND_702;
  reg [31:0] _RAND_703;
  reg [31:0] _RAND_704;
  reg [31:0] _RAND_705;
  reg [31:0] _RAND_706;
  reg [31:0] _RAND_707;
  reg [31:0] _RAND_708;
  reg [31:0] _RAND_709;
  reg [31:0] _RAND_710;
  reg [31:0] _RAND_711;
  reg [31:0] _RAND_712;
  reg [31:0] _RAND_713;
  reg [31:0] _RAND_714;
  reg [31:0] _RAND_715;
  reg [31:0] _RAND_716;
  reg [31:0] _RAND_717;
  reg [31:0] _RAND_718;
  reg [31:0] _RAND_719;
  reg [31:0] _RAND_720;
  reg [31:0] _RAND_721;
  reg [31:0] _RAND_722;
  reg [31:0] _RAND_723;
  reg [31:0] _RAND_724;
  reg [31:0] _RAND_725;
  reg [31:0] _RAND_726;
  reg [31:0] _RAND_727;
  reg [31:0] _RAND_728;
  reg [31:0] _RAND_729;
  reg [31:0] _RAND_730;
  reg [31:0] _RAND_731;
  reg [31:0] _RAND_732;
  reg [31:0] _RAND_733;
  reg [31:0] _RAND_734;
  reg [31:0] _RAND_735;
  reg [31:0] _RAND_736;
  reg [31:0] _RAND_737;
  reg [31:0] _RAND_738;
  reg [31:0] _RAND_739;
  reg [31:0] _RAND_740;
  reg [31:0] _RAND_741;
  reg [31:0] _RAND_742;
  reg [31:0] _RAND_743;
  reg [31:0] _RAND_744;
  reg [31:0] _RAND_745;
  reg [31:0] _RAND_746;
  reg [31:0] _RAND_747;
  reg [31:0] _RAND_748;
  reg [31:0] _RAND_749;
  reg [31:0] _RAND_750;
  reg [31:0] _RAND_751;
  reg [31:0] _RAND_752;
  reg [31:0] _RAND_753;
  reg [31:0] _RAND_754;
  reg [31:0] _RAND_755;
  reg [31:0] _RAND_756;
  reg [31:0] _RAND_757;
  reg [31:0] _RAND_758;
  reg [31:0] _RAND_759;
  reg [31:0] _RAND_760;
  reg [31:0] _RAND_761;
  reg [31:0] _RAND_762;
  reg [31:0] _RAND_763;
  reg [31:0] _RAND_764;
  reg [31:0] _RAND_765;
  reg [31:0] _RAND_766;
  reg [31:0] _RAND_767;
  reg [31:0] _RAND_768;
  reg [31:0] _RAND_769;
  reg [31:0] _RAND_770;
  reg [31:0] _RAND_771;
  reg [31:0] _RAND_772;
  reg [31:0] _RAND_773;
  reg [31:0] _RAND_774;
  reg [31:0] _RAND_775;
  reg [31:0] _RAND_776;
  reg [31:0] _RAND_777;
  reg [31:0] _RAND_778;
  reg [31:0] _RAND_779;
  reg [31:0] _RAND_780;
  reg [31:0] _RAND_781;
  reg [31:0] _RAND_782;
  reg [31:0] _RAND_783;
  reg [31:0] _RAND_784;
  reg [31:0] _RAND_785;
  reg [31:0] _RAND_786;
  reg [31:0] _RAND_787;
  reg [31:0] _RAND_788;
  reg [31:0] _RAND_789;
  reg [31:0] _RAND_790;
  reg [31:0] _RAND_791;
  reg [31:0] _RAND_792;
  reg [31:0] _RAND_793;
  reg [31:0] _RAND_794;
  reg [31:0] _RAND_795;
  reg [31:0] _RAND_796;
  reg [31:0] _RAND_797;
  reg [31:0] _RAND_798;
  reg [31:0] _RAND_799;
  reg [31:0] _RAND_800;
  reg [31:0] _RAND_801;
  reg [31:0] _RAND_802;
  reg [31:0] _RAND_803;
  reg [31:0] _RAND_804;
  reg [31:0] _RAND_805;
  reg [31:0] _RAND_806;
  reg [31:0] _RAND_807;
  reg [31:0] _RAND_808;
  reg [31:0] _RAND_809;
  reg [31:0] _RAND_810;
  reg [31:0] _RAND_811;
  reg [31:0] _RAND_812;
  reg [31:0] _RAND_813;
  reg [31:0] _RAND_814;
  reg [31:0] _RAND_815;
  reg [31:0] _RAND_816;
  reg [31:0] _RAND_817;
  reg [31:0] _RAND_818;
  reg [31:0] _RAND_819;
  reg [31:0] _RAND_820;
  reg [31:0] _RAND_821;
  reg [31:0] _RAND_822;
  reg [31:0] _RAND_823;
  reg [31:0] _RAND_824;
  reg [31:0] _RAND_825;
  reg [31:0] _RAND_826;
  reg [31:0] _RAND_827;
  reg [31:0] _RAND_828;
  reg [31:0] _RAND_829;
  reg [31:0] _RAND_830;
  reg [31:0] _RAND_831;
  reg [31:0] _RAND_832;
  reg [31:0] _RAND_833;
  reg [31:0] _RAND_834;
  reg [31:0] _RAND_835;
  reg [31:0] _RAND_836;
  reg [31:0] _RAND_837;
  reg [31:0] _RAND_838;
  reg [31:0] _RAND_839;
  reg [31:0] _RAND_840;
  reg [31:0] _RAND_841;
  reg [31:0] _RAND_842;
  reg [31:0] _RAND_843;
  reg [31:0] _RAND_844;
  reg [31:0] _RAND_845;
  reg [31:0] _RAND_846;
  reg [31:0] _RAND_847;
  reg [31:0] _RAND_848;
  reg [31:0] _RAND_849;
  reg [31:0] _RAND_850;
  reg [31:0] _RAND_851;
  reg [31:0] _RAND_852;
  reg [31:0] _RAND_853;
  reg [31:0] _RAND_854;
  reg [31:0] _RAND_855;
  reg [31:0] _RAND_856;
  reg [31:0] _RAND_857;
  reg [31:0] _RAND_858;
  reg [31:0] _RAND_859;
  reg [31:0] _RAND_860;
  reg [31:0] _RAND_861;
  reg [31:0] _RAND_862;
  reg [31:0] _RAND_863;
  reg [31:0] _RAND_864;
  reg [31:0] _RAND_865;
  reg [31:0] _RAND_866;
  reg [31:0] _RAND_867;
  reg [31:0] _RAND_868;
  reg [31:0] _RAND_869;
  reg [31:0] _RAND_870;
  reg [31:0] _RAND_871;
  reg [31:0] _RAND_872;
  reg [31:0] _RAND_873;
  reg [31:0] _RAND_874;
  reg [31:0] _RAND_875;
  reg [31:0] _RAND_876;
  reg [31:0] _RAND_877;
  reg [31:0] _RAND_878;
  reg [31:0] _RAND_879;
  reg [31:0] _RAND_880;
  reg [31:0] _RAND_881;
  reg [31:0] _RAND_882;
  reg [31:0] _RAND_883;
  reg [31:0] _RAND_884;
  reg [31:0] _RAND_885;
  reg [31:0] _RAND_886;
  reg [31:0] _RAND_887;
  reg [31:0] _RAND_888;
  reg [31:0] _RAND_889;
  reg [31:0] _RAND_890;
  reg [31:0] _RAND_891;
  reg [31:0] _RAND_892;
  reg [31:0] _RAND_893;
  reg [31:0] _RAND_894;
  reg [31:0] _RAND_895;
  reg [31:0] _RAND_896;
  reg [31:0] _RAND_897;
`endif // RANDOMIZE_REG_INIT
  wire  rs1x0 = io_rs1Addr == 5'h0; // @[bht.scala 45:29]
  wire  rs1x1 = io_rs1Addr == 5'h1; // @[bht.scala 46:29]
  wire [63:0] _rs1x1Data_T_2 = io_wbRdEn & io_wbRdAddr == 5'h1 ? io_wbRdData : io_rs1x1Data; // @[bht.scala 50:28]
  wire [63:0] _rs1x1Data_T_3 = io_memX1En ? io_memAluRes : _rs1x1Data_T_2; // @[bht.scala 49:26]
  wire [63:0] rs1x1Data = io_exeX1En ? io_exeAluRes : _rs1x1Data_T_3; // @[bht.scala 48:24]
  wire [63:0] _op1_T_3 = io_jalr & rs1x1 ? rs1x1Data : io_rs1Data; // @[bht.scala 54:22]
  wire [63:0] _op1_T_4 = io_jalr & rs1x0 ? 64'h0 : _op1_T_3; // @[bht.scala 53:20]
  wire [63:0] op1 = io_bxx | io_jal ? {{32'd0}, io_pc} : _op1_T_4; // @[bht.scala 52:18]
  reg [6:0] ghr; // @[bht.scala 107:22]
  reg [6:0] bht_0; // @[bht.scala 108:22]
  reg [6:0] bht_1; // @[bht.scala 108:22]
  reg [6:0] bht_2; // @[bht.scala 108:22]
  reg [6:0] bht_3; // @[bht.scala 108:22]
  reg [6:0] bht_4; // @[bht.scala 108:22]
  reg [6:0] bht_5; // @[bht.scala 108:22]
  reg [6:0] bht_6; // @[bht.scala 108:22]
  reg [6:0] bht_7; // @[bht.scala 108:22]
  reg [6:0] bht_8; // @[bht.scala 108:22]
  reg [6:0] bht_9; // @[bht.scala 108:22]
  reg [6:0] bht_10; // @[bht.scala 108:22]
  reg [6:0] bht_11; // @[bht.scala 108:22]
  reg [6:0] bht_12; // @[bht.scala 108:22]
  reg [6:0] bht_13; // @[bht.scala 108:22]
  reg [6:0] bht_14; // @[bht.scala 108:22]
  reg [6:0] bht_15; // @[bht.scala 108:22]
  reg [6:0] bht_16; // @[bht.scala 108:22]
  reg [6:0] bht_17; // @[bht.scala 108:22]
  reg [6:0] bht_18; // @[bht.scala 108:22]
  reg [6:0] bht_19; // @[bht.scala 108:22]
  reg [6:0] bht_20; // @[bht.scala 108:22]
  reg [6:0] bht_21; // @[bht.scala 108:22]
  reg [6:0] bht_22; // @[bht.scala 108:22]
  reg [6:0] bht_23; // @[bht.scala 108:22]
  reg [6:0] bht_24; // @[bht.scala 108:22]
  reg [6:0] bht_25; // @[bht.scala 108:22]
  reg [6:0] bht_26; // @[bht.scala 108:22]
  reg [6:0] bht_27; // @[bht.scala 108:22]
  reg [6:0] bht_28; // @[bht.scala 108:22]
  reg [6:0] bht_29; // @[bht.scala 108:22]
  reg [6:0] bht_30; // @[bht.scala 108:22]
  reg [6:0] bht_31; // @[bht.scala 108:22]
  reg [6:0] bht_32; // @[bht.scala 108:22]
  reg [6:0] bht_33; // @[bht.scala 108:22]
  reg [6:0] bht_34; // @[bht.scala 108:22]
  reg [6:0] bht_35; // @[bht.scala 108:22]
  reg [6:0] bht_36; // @[bht.scala 108:22]
  reg [6:0] bht_37; // @[bht.scala 108:22]
  reg [6:0] bht_38; // @[bht.scala 108:22]
  reg [6:0] bht_39; // @[bht.scala 108:22]
  reg [6:0] bht_40; // @[bht.scala 108:22]
  reg [6:0] bht_41; // @[bht.scala 108:22]
  reg [6:0] bht_42; // @[bht.scala 108:22]
  reg [6:0] bht_43; // @[bht.scala 108:22]
  reg [6:0] bht_44; // @[bht.scala 108:22]
  reg [6:0] bht_45; // @[bht.scala 108:22]
  reg [6:0] bht_46; // @[bht.scala 108:22]
  reg [6:0] bht_47; // @[bht.scala 108:22]
  reg [6:0] bht_48; // @[bht.scala 108:22]
  reg [6:0] bht_49; // @[bht.scala 108:22]
  reg [6:0] bht_50; // @[bht.scala 108:22]
  reg [6:0] bht_51; // @[bht.scala 108:22]
  reg [6:0] bht_52; // @[bht.scala 108:22]
  reg [6:0] bht_53; // @[bht.scala 108:22]
  reg [6:0] bht_54; // @[bht.scala 108:22]
  reg [6:0] bht_55; // @[bht.scala 108:22]
  reg [6:0] bht_56; // @[bht.scala 108:22]
  reg [6:0] bht_57; // @[bht.scala 108:22]
  reg [6:0] bht_58; // @[bht.scala 108:22]
  reg [6:0] bht_59; // @[bht.scala 108:22]
  reg [6:0] bht_60; // @[bht.scala 108:22]
  reg [6:0] bht_61; // @[bht.scala 108:22]
  reg [6:0] bht_62; // @[bht.scala 108:22]
  reg [6:0] bht_63; // @[bht.scala 108:22]
  reg [6:0] bht_64; // @[bht.scala 108:22]
  reg [6:0] bht_65; // @[bht.scala 108:22]
  reg [6:0] bht_66; // @[bht.scala 108:22]
  reg [6:0] bht_67; // @[bht.scala 108:22]
  reg [6:0] bht_68; // @[bht.scala 108:22]
  reg [6:0] bht_69; // @[bht.scala 108:22]
  reg [6:0] bht_70; // @[bht.scala 108:22]
  reg [6:0] bht_71; // @[bht.scala 108:22]
  reg [6:0] bht_72; // @[bht.scala 108:22]
  reg [6:0] bht_73; // @[bht.scala 108:22]
  reg [6:0] bht_74; // @[bht.scala 108:22]
  reg [6:0] bht_75; // @[bht.scala 108:22]
  reg [6:0] bht_76; // @[bht.scala 108:22]
  reg [6:0] bht_77; // @[bht.scala 108:22]
  reg [6:0] bht_78; // @[bht.scala 108:22]
  reg [6:0] bht_79; // @[bht.scala 108:22]
  reg [6:0] bht_80; // @[bht.scala 108:22]
  reg [6:0] bht_81; // @[bht.scala 108:22]
  reg [6:0] bht_82; // @[bht.scala 108:22]
  reg [6:0] bht_83; // @[bht.scala 108:22]
  reg [6:0] bht_84; // @[bht.scala 108:22]
  reg [6:0] bht_85; // @[bht.scala 108:22]
  reg [6:0] bht_86; // @[bht.scala 108:22]
  reg [6:0] bht_87; // @[bht.scala 108:22]
  reg [6:0] bht_88; // @[bht.scala 108:22]
  reg [6:0] bht_89; // @[bht.scala 108:22]
  reg [6:0] bht_90; // @[bht.scala 108:22]
  reg [6:0] bht_91; // @[bht.scala 108:22]
  reg [6:0] bht_92; // @[bht.scala 108:22]
  reg [6:0] bht_93; // @[bht.scala 108:22]
  reg [6:0] bht_94; // @[bht.scala 108:22]
  reg [6:0] bht_95; // @[bht.scala 108:22]
  reg [6:0] bht_96; // @[bht.scala 108:22]
  reg [6:0] bht_97; // @[bht.scala 108:22]
  reg [6:0] bht_98; // @[bht.scala 108:22]
  reg [6:0] bht_99; // @[bht.scala 108:22]
  reg [6:0] bht_100; // @[bht.scala 108:22]
  reg [6:0] bht_101; // @[bht.scala 108:22]
  reg [6:0] bht_102; // @[bht.scala 108:22]
  reg [6:0] bht_103; // @[bht.scala 108:22]
  reg [6:0] bht_104; // @[bht.scala 108:22]
  reg [6:0] bht_105; // @[bht.scala 108:22]
  reg [6:0] bht_106; // @[bht.scala 108:22]
  reg [6:0] bht_107; // @[bht.scala 108:22]
  reg [6:0] bht_108; // @[bht.scala 108:22]
  reg [6:0] bht_109; // @[bht.scala 108:22]
  reg [6:0] bht_110; // @[bht.scala 108:22]
  reg [6:0] bht_111; // @[bht.scala 108:22]
  reg [6:0] bht_112; // @[bht.scala 108:22]
  reg [6:0] bht_113; // @[bht.scala 108:22]
  reg [6:0] bht_114; // @[bht.scala 108:22]
  reg [6:0] bht_115; // @[bht.scala 108:22]
  reg [6:0] bht_116; // @[bht.scala 108:22]
  reg [6:0] bht_117; // @[bht.scala 108:22]
  reg [6:0] bht_118; // @[bht.scala 108:22]
  reg [6:0] bht_119; // @[bht.scala 108:22]
  reg [6:0] bht_120; // @[bht.scala 108:22]
  reg [6:0] bht_121; // @[bht.scala 108:22]
  reg [6:0] bht_122; // @[bht.scala 108:22]
  reg [6:0] bht_123; // @[bht.scala 108:22]
  reg [6:0] bht_124; // @[bht.scala 108:22]
  reg [6:0] bht_125; // @[bht.scala 108:22]
  reg [6:0] bht_126; // @[bht.scala 108:22]
  reg [6:0] bht_127; // @[bht.scala 108:22]
  reg [1:0] pht_0_0; // @[bht.scala 109:22]
  reg [1:0] pht_0_1; // @[bht.scala 109:22]
  reg [1:0] pht_0_2; // @[bht.scala 109:22]
  reg [1:0] pht_0_3; // @[bht.scala 109:22]
  reg [1:0] pht_0_4; // @[bht.scala 109:22]
  reg [1:0] pht_0_5; // @[bht.scala 109:22]
  reg [1:0] pht_0_6; // @[bht.scala 109:22]
  reg [1:0] pht_0_7; // @[bht.scala 109:22]
  reg [1:0] pht_0_8; // @[bht.scala 109:22]
  reg [1:0] pht_0_9; // @[bht.scala 109:22]
  reg [1:0] pht_0_10; // @[bht.scala 109:22]
  reg [1:0] pht_0_11; // @[bht.scala 109:22]
  reg [1:0] pht_0_12; // @[bht.scala 109:22]
  reg [1:0] pht_0_13; // @[bht.scala 109:22]
  reg [1:0] pht_0_14; // @[bht.scala 109:22]
  reg [1:0] pht_0_15; // @[bht.scala 109:22]
  reg [1:0] pht_0_16; // @[bht.scala 109:22]
  reg [1:0] pht_0_17; // @[bht.scala 109:22]
  reg [1:0] pht_0_18; // @[bht.scala 109:22]
  reg [1:0] pht_0_19; // @[bht.scala 109:22]
  reg [1:0] pht_0_20; // @[bht.scala 109:22]
  reg [1:0] pht_0_21; // @[bht.scala 109:22]
  reg [1:0] pht_0_22; // @[bht.scala 109:22]
  reg [1:0] pht_0_23; // @[bht.scala 109:22]
  reg [1:0] pht_0_24; // @[bht.scala 109:22]
  reg [1:0] pht_0_25; // @[bht.scala 109:22]
  reg [1:0] pht_0_26; // @[bht.scala 109:22]
  reg [1:0] pht_0_27; // @[bht.scala 109:22]
  reg [1:0] pht_0_28; // @[bht.scala 109:22]
  reg [1:0] pht_0_29; // @[bht.scala 109:22]
  reg [1:0] pht_0_30; // @[bht.scala 109:22]
  reg [1:0] pht_0_31; // @[bht.scala 109:22]
  reg [1:0] pht_0_32; // @[bht.scala 109:22]
  reg [1:0] pht_0_33; // @[bht.scala 109:22]
  reg [1:0] pht_0_34; // @[bht.scala 109:22]
  reg [1:0] pht_0_35; // @[bht.scala 109:22]
  reg [1:0] pht_0_36; // @[bht.scala 109:22]
  reg [1:0] pht_0_37; // @[bht.scala 109:22]
  reg [1:0] pht_0_38; // @[bht.scala 109:22]
  reg [1:0] pht_0_39; // @[bht.scala 109:22]
  reg [1:0] pht_0_40; // @[bht.scala 109:22]
  reg [1:0] pht_0_41; // @[bht.scala 109:22]
  reg [1:0] pht_0_42; // @[bht.scala 109:22]
  reg [1:0] pht_0_43; // @[bht.scala 109:22]
  reg [1:0] pht_0_44; // @[bht.scala 109:22]
  reg [1:0] pht_0_45; // @[bht.scala 109:22]
  reg [1:0] pht_0_46; // @[bht.scala 109:22]
  reg [1:0] pht_0_47; // @[bht.scala 109:22]
  reg [1:0] pht_0_48; // @[bht.scala 109:22]
  reg [1:0] pht_0_49; // @[bht.scala 109:22]
  reg [1:0] pht_0_50; // @[bht.scala 109:22]
  reg [1:0] pht_0_51; // @[bht.scala 109:22]
  reg [1:0] pht_0_52; // @[bht.scala 109:22]
  reg [1:0] pht_0_53; // @[bht.scala 109:22]
  reg [1:0] pht_0_54; // @[bht.scala 109:22]
  reg [1:0] pht_0_55; // @[bht.scala 109:22]
  reg [1:0] pht_0_56; // @[bht.scala 109:22]
  reg [1:0] pht_0_57; // @[bht.scala 109:22]
  reg [1:0] pht_0_58; // @[bht.scala 109:22]
  reg [1:0] pht_0_59; // @[bht.scala 109:22]
  reg [1:0] pht_0_60; // @[bht.scala 109:22]
  reg [1:0] pht_0_61; // @[bht.scala 109:22]
  reg [1:0] pht_0_62; // @[bht.scala 109:22]
  reg [1:0] pht_0_63; // @[bht.scala 109:22]
  reg [1:0] pht_0_64; // @[bht.scala 109:22]
  reg [1:0] pht_0_65; // @[bht.scala 109:22]
  reg [1:0] pht_0_66; // @[bht.scala 109:22]
  reg [1:0] pht_0_67; // @[bht.scala 109:22]
  reg [1:0] pht_0_68; // @[bht.scala 109:22]
  reg [1:0] pht_0_69; // @[bht.scala 109:22]
  reg [1:0] pht_0_70; // @[bht.scala 109:22]
  reg [1:0] pht_0_71; // @[bht.scala 109:22]
  reg [1:0] pht_0_72; // @[bht.scala 109:22]
  reg [1:0] pht_0_73; // @[bht.scala 109:22]
  reg [1:0] pht_0_74; // @[bht.scala 109:22]
  reg [1:0] pht_0_75; // @[bht.scala 109:22]
  reg [1:0] pht_0_76; // @[bht.scala 109:22]
  reg [1:0] pht_0_77; // @[bht.scala 109:22]
  reg [1:0] pht_0_78; // @[bht.scala 109:22]
  reg [1:0] pht_0_79; // @[bht.scala 109:22]
  reg [1:0] pht_0_80; // @[bht.scala 109:22]
  reg [1:0] pht_0_81; // @[bht.scala 109:22]
  reg [1:0] pht_0_82; // @[bht.scala 109:22]
  reg [1:0] pht_0_83; // @[bht.scala 109:22]
  reg [1:0] pht_0_84; // @[bht.scala 109:22]
  reg [1:0] pht_0_85; // @[bht.scala 109:22]
  reg [1:0] pht_0_86; // @[bht.scala 109:22]
  reg [1:0] pht_0_87; // @[bht.scala 109:22]
  reg [1:0] pht_0_88; // @[bht.scala 109:22]
  reg [1:0] pht_0_89; // @[bht.scala 109:22]
  reg [1:0] pht_0_90; // @[bht.scala 109:22]
  reg [1:0] pht_0_91; // @[bht.scala 109:22]
  reg [1:0] pht_0_92; // @[bht.scala 109:22]
  reg [1:0] pht_0_93; // @[bht.scala 109:22]
  reg [1:0] pht_0_94; // @[bht.scala 109:22]
  reg [1:0] pht_0_95; // @[bht.scala 109:22]
  reg [1:0] pht_0_96; // @[bht.scala 109:22]
  reg [1:0] pht_0_97; // @[bht.scala 109:22]
  reg [1:0] pht_0_98; // @[bht.scala 109:22]
  reg [1:0] pht_0_99; // @[bht.scala 109:22]
  reg [1:0] pht_0_100; // @[bht.scala 109:22]
  reg [1:0] pht_0_101; // @[bht.scala 109:22]
  reg [1:0] pht_0_102; // @[bht.scala 109:22]
  reg [1:0] pht_0_103; // @[bht.scala 109:22]
  reg [1:0] pht_0_104; // @[bht.scala 109:22]
  reg [1:0] pht_0_105; // @[bht.scala 109:22]
  reg [1:0] pht_0_106; // @[bht.scala 109:22]
  reg [1:0] pht_0_107; // @[bht.scala 109:22]
  reg [1:0] pht_0_108; // @[bht.scala 109:22]
  reg [1:0] pht_0_109; // @[bht.scala 109:22]
  reg [1:0] pht_0_110; // @[bht.scala 109:22]
  reg [1:0] pht_0_111; // @[bht.scala 109:22]
  reg [1:0] pht_0_112; // @[bht.scala 109:22]
  reg [1:0] pht_0_113; // @[bht.scala 109:22]
  reg [1:0] pht_0_114; // @[bht.scala 109:22]
  reg [1:0] pht_0_115; // @[bht.scala 109:22]
  reg [1:0] pht_0_116; // @[bht.scala 109:22]
  reg [1:0] pht_0_117; // @[bht.scala 109:22]
  reg [1:0] pht_0_118; // @[bht.scala 109:22]
  reg [1:0] pht_0_119; // @[bht.scala 109:22]
  reg [1:0] pht_0_120; // @[bht.scala 109:22]
  reg [1:0] pht_0_121; // @[bht.scala 109:22]
  reg [1:0] pht_0_122; // @[bht.scala 109:22]
  reg [1:0] pht_0_123; // @[bht.scala 109:22]
  reg [1:0] pht_0_124; // @[bht.scala 109:22]
  reg [1:0] pht_0_125; // @[bht.scala 109:22]
  reg [1:0] pht_0_126; // @[bht.scala 109:22]
  reg [1:0] pht_0_127; // @[bht.scala 109:22]
  reg [1:0] pht_1_0; // @[bht.scala 109:22]
  reg [1:0] pht_1_1; // @[bht.scala 109:22]
  reg [1:0] pht_1_2; // @[bht.scala 109:22]
  reg [1:0] pht_1_3; // @[bht.scala 109:22]
  reg [1:0] pht_1_4; // @[bht.scala 109:22]
  reg [1:0] pht_1_5; // @[bht.scala 109:22]
  reg [1:0] pht_1_6; // @[bht.scala 109:22]
  reg [1:0] pht_1_7; // @[bht.scala 109:22]
  reg [1:0] pht_1_8; // @[bht.scala 109:22]
  reg [1:0] pht_1_9; // @[bht.scala 109:22]
  reg [1:0] pht_1_10; // @[bht.scala 109:22]
  reg [1:0] pht_1_11; // @[bht.scala 109:22]
  reg [1:0] pht_1_12; // @[bht.scala 109:22]
  reg [1:0] pht_1_13; // @[bht.scala 109:22]
  reg [1:0] pht_1_14; // @[bht.scala 109:22]
  reg [1:0] pht_1_15; // @[bht.scala 109:22]
  reg [1:0] pht_1_16; // @[bht.scala 109:22]
  reg [1:0] pht_1_17; // @[bht.scala 109:22]
  reg [1:0] pht_1_18; // @[bht.scala 109:22]
  reg [1:0] pht_1_19; // @[bht.scala 109:22]
  reg [1:0] pht_1_20; // @[bht.scala 109:22]
  reg [1:0] pht_1_21; // @[bht.scala 109:22]
  reg [1:0] pht_1_22; // @[bht.scala 109:22]
  reg [1:0] pht_1_23; // @[bht.scala 109:22]
  reg [1:0] pht_1_24; // @[bht.scala 109:22]
  reg [1:0] pht_1_25; // @[bht.scala 109:22]
  reg [1:0] pht_1_26; // @[bht.scala 109:22]
  reg [1:0] pht_1_27; // @[bht.scala 109:22]
  reg [1:0] pht_1_28; // @[bht.scala 109:22]
  reg [1:0] pht_1_29; // @[bht.scala 109:22]
  reg [1:0] pht_1_30; // @[bht.scala 109:22]
  reg [1:0] pht_1_31; // @[bht.scala 109:22]
  reg [1:0] pht_1_32; // @[bht.scala 109:22]
  reg [1:0] pht_1_33; // @[bht.scala 109:22]
  reg [1:0] pht_1_34; // @[bht.scala 109:22]
  reg [1:0] pht_1_35; // @[bht.scala 109:22]
  reg [1:0] pht_1_36; // @[bht.scala 109:22]
  reg [1:0] pht_1_37; // @[bht.scala 109:22]
  reg [1:0] pht_1_38; // @[bht.scala 109:22]
  reg [1:0] pht_1_39; // @[bht.scala 109:22]
  reg [1:0] pht_1_40; // @[bht.scala 109:22]
  reg [1:0] pht_1_41; // @[bht.scala 109:22]
  reg [1:0] pht_1_42; // @[bht.scala 109:22]
  reg [1:0] pht_1_43; // @[bht.scala 109:22]
  reg [1:0] pht_1_44; // @[bht.scala 109:22]
  reg [1:0] pht_1_45; // @[bht.scala 109:22]
  reg [1:0] pht_1_46; // @[bht.scala 109:22]
  reg [1:0] pht_1_47; // @[bht.scala 109:22]
  reg [1:0] pht_1_48; // @[bht.scala 109:22]
  reg [1:0] pht_1_49; // @[bht.scala 109:22]
  reg [1:0] pht_1_50; // @[bht.scala 109:22]
  reg [1:0] pht_1_51; // @[bht.scala 109:22]
  reg [1:0] pht_1_52; // @[bht.scala 109:22]
  reg [1:0] pht_1_53; // @[bht.scala 109:22]
  reg [1:0] pht_1_54; // @[bht.scala 109:22]
  reg [1:0] pht_1_55; // @[bht.scala 109:22]
  reg [1:0] pht_1_56; // @[bht.scala 109:22]
  reg [1:0] pht_1_57; // @[bht.scala 109:22]
  reg [1:0] pht_1_58; // @[bht.scala 109:22]
  reg [1:0] pht_1_59; // @[bht.scala 109:22]
  reg [1:0] pht_1_60; // @[bht.scala 109:22]
  reg [1:0] pht_1_61; // @[bht.scala 109:22]
  reg [1:0] pht_1_62; // @[bht.scala 109:22]
  reg [1:0] pht_1_63; // @[bht.scala 109:22]
  reg [1:0] pht_1_64; // @[bht.scala 109:22]
  reg [1:0] pht_1_65; // @[bht.scala 109:22]
  reg [1:0] pht_1_66; // @[bht.scala 109:22]
  reg [1:0] pht_1_67; // @[bht.scala 109:22]
  reg [1:0] pht_1_68; // @[bht.scala 109:22]
  reg [1:0] pht_1_69; // @[bht.scala 109:22]
  reg [1:0] pht_1_70; // @[bht.scala 109:22]
  reg [1:0] pht_1_71; // @[bht.scala 109:22]
  reg [1:0] pht_1_72; // @[bht.scala 109:22]
  reg [1:0] pht_1_73; // @[bht.scala 109:22]
  reg [1:0] pht_1_74; // @[bht.scala 109:22]
  reg [1:0] pht_1_75; // @[bht.scala 109:22]
  reg [1:0] pht_1_76; // @[bht.scala 109:22]
  reg [1:0] pht_1_77; // @[bht.scala 109:22]
  reg [1:0] pht_1_78; // @[bht.scala 109:22]
  reg [1:0] pht_1_79; // @[bht.scala 109:22]
  reg [1:0] pht_1_80; // @[bht.scala 109:22]
  reg [1:0] pht_1_81; // @[bht.scala 109:22]
  reg [1:0] pht_1_82; // @[bht.scala 109:22]
  reg [1:0] pht_1_83; // @[bht.scala 109:22]
  reg [1:0] pht_1_84; // @[bht.scala 109:22]
  reg [1:0] pht_1_85; // @[bht.scala 109:22]
  reg [1:0] pht_1_86; // @[bht.scala 109:22]
  reg [1:0] pht_1_87; // @[bht.scala 109:22]
  reg [1:0] pht_1_88; // @[bht.scala 109:22]
  reg [1:0] pht_1_89; // @[bht.scala 109:22]
  reg [1:0] pht_1_90; // @[bht.scala 109:22]
  reg [1:0] pht_1_91; // @[bht.scala 109:22]
  reg [1:0] pht_1_92; // @[bht.scala 109:22]
  reg [1:0] pht_1_93; // @[bht.scala 109:22]
  reg [1:0] pht_1_94; // @[bht.scala 109:22]
  reg [1:0] pht_1_95; // @[bht.scala 109:22]
  reg [1:0] pht_1_96; // @[bht.scala 109:22]
  reg [1:0] pht_1_97; // @[bht.scala 109:22]
  reg [1:0] pht_1_98; // @[bht.scala 109:22]
  reg [1:0] pht_1_99; // @[bht.scala 109:22]
  reg [1:0] pht_1_100; // @[bht.scala 109:22]
  reg [1:0] pht_1_101; // @[bht.scala 109:22]
  reg [1:0] pht_1_102; // @[bht.scala 109:22]
  reg [1:0] pht_1_103; // @[bht.scala 109:22]
  reg [1:0] pht_1_104; // @[bht.scala 109:22]
  reg [1:0] pht_1_105; // @[bht.scala 109:22]
  reg [1:0] pht_1_106; // @[bht.scala 109:22]
  reg [1:0] pht_1_107; // @[bht.scala 109:22]
  reg [1:0] pht_1_108; // @[bht.scala 109:22]
  reg [1:0] pht_1_109; // @[bht.scala 109:22]
  reg [1:0] pht_1_110; // @[bht.scala 109:22]
  reg [1:0] pht_1_111; // @[bht.scala 109:22]
  reg [1:0] pht_1_112; // @[bht.scala 109:22]
  reg [1:0] pht_1_113; // @[bht.scala 109:22]
  reg [1:0] pht_1_114; // @[bht.scala 109:22]
  reg [1:0] pht_1_115; // @[bht.scala 109:22]
  reg [1:0] pht_1_116; // @[bht.scala 109:22]
  reg [1:0] pht_1_117; // @[bht.scala 109:22]
  reg [1:0] pht_1_118; // @[bht.scala 109:22]
  reg [1:0] pht_1_119; // @[bht.scala 109:22]
  reg [1:0] pht_1_120; // @[bht.scala 109:22]
  reg [1:0] pht_1_121; // @[bht.scala 109:22]
  reg [1:0] pht_1_122; // @[bht.scala 109:22]
  reg [1:0] pht_1_123; // @[bht.scala 109:22]
  reg [1:0] pht_1_124; // @[bht.scala 109:22]
  reg [1:0] pht_1_125; // @[bht.scala 109:22]
  reg [1:0] pht_1_126; // @[bht.scala 109:22]
  reg [1:0] pht_1_127; // @[bht.scala 109:22]
  reg [1:0] pht_2_0; // @[bht.scala 109:22]
  reg [1:0] pht_2_1; // @[bht.scala 109:22]
  reg [1:0] pht_2_2; // @[bht.scala 109:22]
  reg [1:0] pht_2_3; // @[bht.scala 109:22]
  reg [1:0] pht_2_4; // @[bht.scala 109:22]
  reg [1:0] pht_2_5; // @[bht.scala 109:22]
  reg [1:0] pht_2_6; // @[bht.scala 109:22]
  reg [1:0] pht_2_7; // @[bht.scala 109:22]
  reg [1:0] pht_2_8; // @[bht.scala 109:22]
  reg [1:0] pht_2_9; // @[bht.scala 109:22]
  reg [1:0] pht_2_10; // @[bht.scala 109:22]
  reg [1:0] pht_2_11; // @[bht.scala 109:22]
  reg [1:0] pht_2_12; // @[bht.scala 109:22]
  reg [1:0] pht_2_13; // @[bht.scala 109:22]
  reg [1:0] pht_2_14; // @[bht.scala 109:22]
  reg [1:0] pht_2_15; // @[bht.scala 109:22]
  reg [1:0] pht_2_16; // @[bht.scala 109:22]
  reg [1:0] pht_2_17; // @[bht.scala 109:22]
  reg [1:0] pht_2_18; // @[bht.scala 109:22]
  reg [1:0] pht_2_19; // @[bht.scala 109:22]
  reg [1:0] pht_2_20; // @[bht.scala 109:22]
  reg [1:0] pht_2_21; // @[bht.scala 109:22]
  reg [1:0] pht_2_22; // @[bht.scala 109:22]
  reg [1:0] pht_2_23; // @[bht.scala 109:22]
  reg [1:0] pht_2_24; // @[bht.scala 109:22]
  reg [1:0] pht_2_25; // @[bht.scala 109:22]
  reg [1:0] pht_2_26; // @[bht.scala 109:22]
  reg [1:0] pht_2_27; // @[bht.scala 109:22]
  reg [1:0] pht_2_28; // @[bht.scala 109:22]
  reg [1:0] pht_2_29; // @[bht.scala 109:22]
  reg [1:0] pht_2_30; // @[bht.scala 109:22]
  reg [1:0] pht_2_31; // @[bht.scala 109:22]
  reg [1:0] pht_2_32; // @[bht.scala 109:22]
  reg [1:0] pht_2_33; // @[bht.scala 109:22]
  reg [1:0] pht_2_34; // @[bht.scala 109:22]
  reg [1:0] pht_2_35; // @[bht.scala 109:22]
  reg [1:0] pht_2_36; // @[bht.scala 109:22]
  reg [1:0] pht_2_37; // @[bht.scala 109:22]
  reg [1:0] pht_2_38; // @[bht.scala 109:22]
  reg [1:0] pht_2_39; // @[bht.scala 109:22]
  reg [1:0] pht_2_40; // @[bht.scala 109:22]
  reg [1:0] pht_2_41; // @[bht.scala 109:22]
  reg [1:0] pht_2_42; // @[bht.scala 109:22]
  reg [1:0] pht_2_43; // @[bht.scala 109:22]
  reg [1:0] pht_2_44; // @[bht.scala 109:22]
  reg [1:0] pht_2_45; // @[bht.scala 109:22]
  reg [1:0] pht_2_46; // @[bht.scala 109:22]
  reg [1:0] pht_2_47; // @[bht.scala 109:22]
  reg [1:0] pht_2_48; // @[bht.scala 109:22]
  reg [1:0] pht_2_49; // @[bht.scala 109:22]
  reg [1:0] pht_2_50; // @[bht.scala 109:22]
  reg [1:0] pht_2_51; // @[bht.scala 109:22]
  reg [1:0] pht_2_52; // @[bht.scala 109:22]
  reg [1:0] pht_2_53; // @[bht.scala 109:22]
  reg [1:0] pht_2_54; // @[bht.scala 109:22]
  reg [1:0] pht_2_55; // @[bht.scala 109:22]
  reg [1:0] pht_2_56; // @[bht.scala 109:22]
  reg [1:0] pht_2_57; // @[bht.scala 109:22]
  reg [1:0] pht_2_58; // @[bht.scala 109:22]
  reg [1:0] pht_2_59; // @[bht.scala 109:22]
  reg [1:0] pht_2_60; // @[bht.scala 109:22]
  reg [1:0] pht_2_61; // @[bht.scala 109:22]
  reg [1:0] pht_2_62; // @[bht.scala 109:22]
  reg [1:0] pht_2_63; // @[bht.scala 109:22]
  reg [1:0] pht_2_64; // @[bht.scala 109:22]
  reg [1:0] pht_2_65; // @[bht.scala 109:22]
  reg [1:0] pht_2_66; // @[bht.scala 109:22]
  reg [1:0] pht_2_67; // @[bht.scala 109:22]
  reg [1:0] pht_2_68; // @[bht.scala 109:22]
  reg [1:0] pht_2_69; // @[bht.scala 109:22]
  reg [1:0] pht_2_70; // @[bht.scala 109:22]
  reg [1:0] pht_2_71; // @[bht.scala 109:22]
  reg [1:0] pht_2_72; // @[bht.scala 109:22]
  reg [1:0] pht_2_73; // @[bht.scala 109:22]
  reg [1:0] pht_2_74; // @[bht.scala 109:22]
  reg [1:0] pht_2_75; // @[bht.scala 109:22]
  reg [1:0] pht_2_76; // @[bht.scala 109:22]
  reg [1:0] pht_2_77; // @[bht.scala 109:22]
  reg [1:0] pht_2_78; // @[bht.scala 109:22]
  reg [1:0] pht_2_79; // @[bht.scala 109:22]
  reg [1:0] pht_2_80; // @[bht.scala 109:22]
  reg [1:0] pht_2_81; // @[bht.scala 109:22]
  reg [1:0] pht_2_82; // @[bht.scala 109:22]
  reg [1:0] pht_2_83; // @[bht.scala 109:22]
  reg [1:0] pht_2_84; // @[bht.scala 109:22]
  reg [1:0] pht_2_85; // @[bht.scala 109:22]
  reg [1:0] pht_2_86; // @[bht.scala 109:22]
  reg [1:0] pht_2_87; // @[bht.scala 109:22]
  reg [1:0] pht_2_88; // @[bht.scala 109:22]
  reg [1:0] pht_2_89; // @[bht.scala 109:22]
  reg [1:0] pht_2_90; // @[bht.scala 109:22]
  reg [1:0] pht_2_91; // @[bht.scala 109:22]
  reg [1:0] pht_2_92; // @[bht.scala 109:22]
  reg [1:0] pht_2_93; // @[bht.scala 109:22]
  reg [1:0] pht_2_94; // @[bht.scala 109:22]
  reg [1:0] pht_2_95; // @[bht.scala 109:22]
  reg [1:0] pht_2_96; // @[bht.scala 109:22]
  reg [1:0] pht_2_97; // @[bht.scala 109:22]
  reg [1:0] pht_2_98; // @[bht.scala 109:22]
  reg [1:0] pht_2_99; // @[bht.scala 109:22]
  reg [1:0] pht_2_100; // @[bht.scala 109:22]
  reg [1:0] pht_2_101; // @[bht.scala 109:22]
  reg [1:0] pht_2_102; // @[bht.scala 109:22]
  reg [1:0] pht_2_103; // @[bht.scala 109:22]
  reg [1:0] pht_2_104; // @[bht.scala 109:22]
  reg [1:0] pht_2_105; // @[bht.scala 109:22]
  reg [1:0] pht_2_106; // @[bht.scala 109:22]
  reg [1:0] pht_2_107; // @[bht.scala 109:22]
  reg [1:0] pht_2_108; // @[bht.scala 109:22]
  reg [1:0] pht_2_109; // @[bht.scala 109:22]
  reg [1:0] pht_2_110; // @[bht.scala 109:22]
  reg [1:0] pht_2_111; // @[bht.scala 109:22]
  reg [1:0] pht_2_112; // @[bht.scala 109:22]
  reg [1:0] pht_2_113; // @[bht.scala 109:22]
  reg [1:0] pht_2_114; // @[bht.scala 109:22]
  reg [1:0] pht_2_115; // @[bht.scala 109:22]
  reg [1:0] pht_2_116; // @[bht.scala 109:22]
  reg [1:0] pht_2_117; // @[bht.scala 109:22]
  reg [1:0] pht_2_118; // @[bht.scala 109:22]
  reg [1:0] pht_2_119; // @[bht.scala 109:22]
  reg [1:0] pht_2_120; // @[bht.scala 109:22]
  reg [1:0] pht_2_121; // @[bht.scala 109:22]
  reg [1:0] pht_2_122; // @[bht.scala 109:22]
  reg [1:0] pht_2_123; // @[bht.scala 109:22]
  reg [1:0] pht_2_124; // @[bht.scala 109:22]
  reg [1:0] pht_2_125; // @[bht.scala 109:22]
  reg [1:0] pht_2_126; // @[bht.scala 109:22]
  reg [1:0] pht_2_127; // @[bht.scala 109:22]
  reg  btbV_0; // @[bht.scala 112:23]
  reg  btbV_1; // @[bht.scala 112:23]
  reg  btbV_2; // @[bht.scala 112:23]
  reg  btbV_3; // @[bht.scala 112:23]
  reg  btbV_4; // @[bht.scala 112:23]
  reg  btbV_5; // @[bht.scala 112:23]
  reg  btbV_6; // @[bht.scala 112:23]
  reg  btbV_7; // @[bht.scala 112:23]
  reg  btbV_8; // @[bht.scala 112:23]
  reg  btbV_9; // @[bht.scala 112:23]
  reg  btbV_10; // @[bht.scala 112:23]
  reg  btbV_11; // @[bht.scala 112:23]
  reg  btbV_12; // @[bht.scala 112:23]
  reg  btbV_13; // @[bht.scala 112:23]
  reg  btbV_14; // @[bht.scala 112:23]
  reg  btbV_15; // @[bht.scala 112:23]
  reg  btbV_16; // @[bht.scala 112:23]
  reg  btbV_17; // @[bht.scala 112:23]
  reg  btbV_18; // @[bht.scala 112:23]
  reg  btbV_19; // @[bht.scala 112:23]
  reg  btbV_20; // @[bht.scala 112:23]
  reg  btbV_21; // @[bht.scala 112:23]
  reg  btbV_22; // @[bht.scala 112:23]
  reg  btbV_23; // @[bht.scala 112:23]
  reg  btbV_24; // @[bht.scala 112:23]
  reg  btbV_25; // @[bht.scala 112:23]
  reg  btbV_26; // @[bht.scala 112:23]
  reg  btbV_27; // @[bht.scala 112:23]
  reg  btbV_28; // @[bht.scala 112:23]
  reg  btbV_29; // @[bht.scala 112:23]
  reg  btbV_30; // @[bht.scala 112:23]
  reg  btbV_31; // @[bht.scala 112:23]
  reg  btbV_32; // @[bht.scala 112:23]
  reg  btbV_33; // @[bht.scala 112:23]
  reg  btbV_34; // @[bht.scala 112:23]
  reg  btbV_35; // @[bht.scala 112:23]
  reg  btbV_36; // @[bht.scala 112:23]
  reg  btbV_37; // @[bht.scala 112:23]
  reg  btbV_38; // @[bht.scala 112:23]
  reg  btbV_39; // @[bht.scala 112:23]
  reg  btbV_40; // @[bht.scala 112:23]
  reg  btbV_41; // @[bht.scala 112:23]
  reg  btbV_42; // @[bht.scala 112:23]
  reg  btbV_43; // @[bht.scala 112:23]
  reg  btbV_44; // @[bht.scala 112:23]
  reg  btbV_45; // @[bht.scala 112:23]
  reg  btbV_46; // @[bht.scala 112:23]
  reg  btbV_47; // @[bht.scala 112:23]
  reg  btbV_48; // @[bht.scala 112:23]
  reg  btbV_49; // @[bht.scala 112:23]
  reg  btbV_50; // @[bht.scala 112:23]
  reg  btbV_51; // @[bht.scala 112:23]
  reg  btbV_52; // @[bht.scala 112:23]
  reg  btbV_53; // @[bht.scala 112:23]
  reg  btbV_54; // @[bht.scala 112:23]
  reg  btbV_55; // @[bht.scala 112:23]
  reg  btbV_56; // @[bht.scala 112:23]
  reg  btbV_57; // @[bht.scala 112:23]
  reg  btbV_58; // @[bht.scala 112:23]
  reg  btbV_59; // @[bht.scala 112:23]
  reg  btbV_60; // @[bht.scala 112:23]
  reg  btbV_61; // @[bht.scala 112:23]
  reg  btbV_62; // @[bht.scala 112:23]
  reg  btbV_63; // @[bht.scala 112:23]
  reg  btbV_64; // @[bht.scala 112:23]
  reg  btbV_65; // @[bht.scala 112:23]
  reg  btbV_66; // @[bht.scala 112:23]
  reg  btbV_67; // @[bht.scala 112:23]
  reg  btbV_68; // @[bht.scala 112:23]
  reg  btbV_69; // @[bht.scala 112:23]
  reg  btbV_70; // @[bht.scala 112:23]
  reg  btbV_71; // @[bht.scala 112:23]
  reg  btbV_72; // @[bht.scala 112:23]
  reg  btbV_73; // @[bht.scala 112:23]
  reg  btbV_74; // @[bht.scala 112:23]
  reg  btbV_75; // @[bht.scala 112:23]
  reg  btbV_76; // @[bht.scala 112:23]
  reg  btbV_77; // @[bht.scala 112:23]
  reg  btbV_78; // @[bht.scala 112:23]
  reg  btbV_79; // @[bht.scala 112:23]
  reg  btbV_80; // @[bht.scala 112:23]
  reg  btbV_81; // @[bht.scala 112:23]
  reg  btbV_82; // @[bht.scala 112:23]
  reg  btbV_83; // @[bht.scala 112:23]
  reg  btbV_84; // @[bht.scala 112:23]
  reg  btbV_85; // @[bht.scala 112:23]
  reg  btbV_86; // @[bht.scala 112:23]
  reg  btbV_87; // @[bht.scala 112:23]
  reg  btbV_88; // @[bht.scala 112:23]
  reg  btbV_89; // @[bht.scala 112:23]
  reg  btbV_90; // @[bht.scala 112:23]
  reg  btbV_91; // @[bht.scala 112:23]
  reg  btbV_92; // @[bht.scala 112:23]
  reg  btbV_93; // @[bht.scala 112:23]
  reg  btbV_94; // @[bht.scala 112:23]
  reg  btbV_95; // @[bht.scala 112:23]
  reg  btbV_96; // @[bht.scala 112:23]
  reg  btbV_97; // @[bht.scala 112:23]
  reg  btbV_98; // @[bht.scala 112:23]
  reg  btbV_99; // @[bht.scala 112:23]
  reg  btbV_100; // @[bht.scala 112:23]
  reg  btbV_101; // @[bht.scala 112:23]
  reg  btbV_102; // @[bht.scala 112:23]
  reg  btbV_103; // @[bht.scala 112:23]
  reg  btbV_104; // @[bht.scala 112:23]
  reg  btbV_105; // @[bht.scala 112:23]
  reg  btbV_106; // @[bht.scala 112:23]
  reg  btbV_107; // @[bht.scala 112:23]
  reg  btbV_108; // @[bht.scala 112:23]
  reg  btbV_109; // @[bht.scala 112:23]
  reg  btbV_110; // @[bht.scala 112:23]
  reg  btbV_111; // @[bht.scala 112:23]
  reg  btbV_112; // @[bht.scala 112:23]
  reg  btbV_113; // @[bht.scala 112:23]
  reg  btbV_114; // @[bht.scala 112:23]
  reg  btbV_115; // @[bht.scala 112:23]
  reg  btbV_116; // @[bht.scala 112:23]
  reg  btbV_117; // @[bht.scala 112:23]
  reg  btbV_118; // @[bht.scala 112:23]
  reg  btbV_119; // @[bht.scala 112:23]
  reg  btbV_120; // @[bht.scala 112:23]
  reg  btbV_121; // @[bht.scala 112:23]
  reg  btbV_122; // @[bht.scala 112:23]
  reg  btbV_123; // @[bht.scala 112:23]
  reg  btbV_124; // @[bht.scala 112:23]
  reg  btbV_125; // @[bht.scala 112:23]
  reg  btbV_126; // @[bht.scala 112:23]
  reg  btbV_127; // @[bht.scala 112:23]
  reg [6:0] btbTag_0; // @[bht.scala 113:25]
  reg [6:0] btbTag_1; // @[bht.scala 113:25]
  reg [6:0] btbTag_2; // @[bht.scala 113:25]
  reg [6:0] btbTag_3; // @[bht.scala 113:25]
  reg [6:0] btbTag_4; // @[bht.scala 113:25]
  reg [6:0] btbTag_5; // @[bht.scala 113:25]
  reg [6:0] btbTag_6; // @[bht.scala 113:25]
  reg [6:0] btbTag_7; // @[bht.scala 113:25]
  reg [6:0] btbTag_8; // @[bht.scala 113:25]
  reg [6:0] btbTag_9; // @[bht.scala 113:25]
  reg [6:0] btbTag_10; // @[bht.scala 113:25]
  reg [6:0] btbTag_11; // @[bht.scala 113:25]
  reg [6:0] btbTag_12; // @[bht.scala 113:25]
  reg [6:0] btbTag_13; // @[bht.scala 113:25]
  reg [6:0] btbTag_14; // @[bht.scala 113:25]
  reg [6:0] btbTag_15; // @[bht.scala 113:25]
  reg [6:0] btbTag_16; // @[bht.scala 113:25]
  reg [6:0] btbTag_17; // @[bht.scala 113:25]
  reg [6:0] btbTag_18; // @[bht.scala 113:25]
  reg [6:0] btbTag_19; // @[bht.scala 113:25]
  reg [6:0] btbTag_20; // @[bht.scala 113:25]
  reg [6:0] btbTag_21; // @[bht.scala 113:25]
  reg [6:0] btbTag_22; // @[bht.scala 113:25]
  reg [6:0] btbTag_23; // @[bht.scala 113:25]
  reg [6:0] btbTag_24; // @[bht.scala 113:25]
  reg [6:0] btbTag_25; // @[bht.scala 113:25]
  reg [6:0] btbTag_26; // @[bht.scala 113:25]
  reg [6:0] btbTag_27; // @[bht.scala 113:25]
  reg [6:0] btbTag_28; // @[bht.scala 113:25]
  reg [6:0] btbTag_29; // @[bht.scala 113:25]
  reg [6:0] btbTag_30; // @[bht.scala 113:25]
  reg [6:0] btbTag_31; // @[bht.scala 113:25]
  reg [6:0] btbTag_32; // @[bht.scala 113:25]
  reg [6:0] btbTag_33; // @[bht.scala 113:25]
  reg [6:0] btbTag_34; // @[bht.scala 113:25]
  reg [6:0] btbTag_35; // @[bht.scala 113:25]
  reg [6:0] btbTag_36; // @[bht.scala 113:25]
  reg [6:0] btbTag_37; // @[bht.scala 113:25]
  reg [6:0] btbTag_38; // @[bht.scala 113:25]
  reg [6:0] btbTag_39; // @[bht.scala 113:25]
  reg [6:0] btbTag_40; // @[bht.scala 113:25]
  reg [6:0] btbTag_41; // @[bht.scala 113:25]
  reg [6:0] btbTag_42; // @[bht.scala 113:25]
  reg [6:0] btbTag_43; // @[bht.scala 113:25]
  reg [6:0] btbTag_44; // @[bht.scala 113:25]
  reg [6:0] btbTag_45; // @[bht.scala 113:25]
  reg [6:0] btbTag_46; // @[bht.scala 113:25]
  reg [6:0] btbTag_47; // @[bht.scala 113:25]
  reg [6:0] btbTag_48; // @[bht.scala 113:25]
  reg [6:0] btbTag_49; // @[bht.scala 113:25]
  reg [6:0] btbTag_50; // @[bht.scala 113:25]
  reg [6:0] btbTag_51; // @[bht.scala 113:25]
  reg [6:0] btbTag_52; // @[bht.scala 113:25]
  reg [6:0] btbTag_53; // @[bht.scala 113:25]
  reg [6:0] btbTag_54; // @[bht.scala 113:25]
  reg [6:0] btbTag_55; // @[bht.scala 113:25]
  reg [6:0] btbTag_56; // @[bht.scala 113:25]
  reg [6:0] btbTag_57; // @[bht.scala 113:25]
  reg [6:0] btbTag_58; // @[bht.scala 113:25]
  reg [6:0] btbTag_59; // @[bht.scala 113:25]
  reg [6:0] btbTag_60; // @[bht.scala 113:25]
  reg [6:0] btbTag_61; // @[bht.scala 113:25]
  reg [6:0] btbTag_62; // @[bht.scala 113:25]
  reg [6:0] btbTag_63; // @[bht.scala 113:25]
  reg [6:0] btbTag_64; // @[bht.scala 113:25]
  reg [6:0] btbTag_65; // @[bht.scala 113:25]
  reg [6:0] btbTag_66; // @[bht.scala 113:25]
  reg [6:0] btbTag_67; // @[bht.scala 113:25]
  reg [6:0] btbTag_68; // @[bht.scala 113:25]
  reg [6:0] btbTag_69; // @[bht.scala 113:25]
  reg [6:0] btbTag_70; // @[bht.scala 113:25]
  reg [6:0] btbTag_71; // @[bht.scala 113:25]
  reg [6:0] btbTag_72; // @[bht.scala 113:25]
  reg [6:0] btbTag_73; // @[bht.scala 113:25]
  reg [6:0] btbTag_74; // @[bht.scala 113:25]
  reg [6:0] btbTag_75; // @[bht.scala 113:25]
  reg [6:0] btbTag_76; // @[bht.scala 113:25]
  reg [6:0] btbTag_77; // @[bht.scala 113:25]
  reg [6:0] btbTag_78; // @[bht.scala 113:25]
  reg [6:0] btbTag_79; // @[bht.scala 113:25]
  reg [6:0] btbTag_80; // @[bht.scala 113:25]
  reg [6:0] btbTag_81; // @[bht.scala 113:25]
  reg [6:0] btbTag_82; // @[bht.scala 113:25]
  reg [6:0] btbTag_83; // @[bht.scala 113:25]
  reg [6:0] btbTag_84; // @[bht.scala 113:25]
  reg [6:0] btbTag_85; // @[bht.scala 113:25]
  reg [6:0] btbTag_86; // @[bht.scala 113:25]
  reg [6:0] btbTag_87; // @[bht.scala 113:25]
  reg [6:0] btbTag_88; // @[bht.scala 113:25]
  reg [6:0] btbTag_89; // @[bht.scala 113:25]
  reg [6:0] btbTag_90; // @[bht.scala 113:25]
  reg [6:0] btbTag_91; // @[bht.scala 113:25]
  reg [6:0] btbTag_92; // @[bht.scala 113:25]
  reg [6:0] btbTag_93; // @[bht.scala 113:25]
  reg [6:0] btbTag_94; // @[bht.scala 113:25]
  reg [6:0] btbTag_95; // @[bht.scala 113:25]
  reg [6:0] btbTag_96; // @[bht.scala 113:25]
  reg [6:0] btbTag_97; // @[bht.scala 113:25]
  reg [6:0] btbTag_98; // @[bht.scala 113:25]
  reg [6:0] btbTag_99; // @[bht.scala 113:25]
  reg [6:0] btbTag_100; // @[bht.scala 113:25]
  reg [6:0] btbTag_101; // @[bht.scala 113:25]
  reg [6:0] btbTag_102; // @[bht.scala 113:25]
  reg [6:0] btbTag_103; // @[bht.scala 113:25]
  reg [6:0] btbTag_104; // @[bht.scala 113:25]
  reg [6:0] btbTag_105; // @[bht.scala 113:25]
  reg [6:0] btbTag_106; // @[bht.scala 113:25]
  reg [6:0] btbTag_107; // @[bht.scala 113:25]
  reg [6:0] btbTag_108; // @[bht.scala 113:25]
  reg [6:0] btbTag_109; // @[bht.scala 113:25]
  reg [6:0] btbTag_110; // @[bht.scala 113:25]
  reg [6:0] btbTag_111; // @[bht.scala 113:25]
  reg [6:0] btbTag_112; // @[bht.scala 113:25]
  reg [6:0] btbTag_113; // @[bht.scala 113:25]
  reg [6:0] btbTag_114; // @[bht.scala 113:25]
  reg [6:0] btbTag_115; // @[bht.scala 113:25]
  reg [6:0] btbTag_116; // @[bht.scala 113:25]
  reg [6:0] btbTag_117; // @[bht.scala 113:25]
  reg [6:0] btbTag_118; // @[bht.scala 113:25]
  reg [6:0] btbTag_119; // @[bht.scala 113:25]
  reg [6:0] btbTag_120; // @[bht.scala 113:25]
  reg [6:0] btbTag_121; // @[bht.scala 113:25]
  reg [6:0] btbTag_122; // @[bht.scala 113:25]
  reg [6:0] btbTag_123; // @[bht.scala 113:25]
  reg [6:0] btbTag_124; // @[bht.scala 113:25]
  reg [6:0] btbTag_125; // @[bht.scala 113:25]
  reg [6:0] btbTag_126; // @[bht.scala 113:25]
  reg [6:0] btbTag_127; // @[bht.scala 113:25]
  reg [31:0] btbMeta_0; // @[bht.scala 114:26]
  reg [31:0] btbMeta_1; // @[bht.scala 114:26]
  reg [31:0] btbMeta_2; // @[bht.scala 114:26]
  reg [31:0] btbMeta_3; // @[bht.scala 114:26]
  reg [31:0] btbMeta_4; // @[bht.scala 114:26]
  reg [31:0] btbMeta_5; // @[bht.scala 114:26]
  reg [31:0] btbMeta_6; // @[bht.scala 114:26]
  reg [31:0] btbMeta_7; // @[bht.scala 114:26]
  reg [31:0] btbMeta_8; // @[bht.scala 114:26]
  reg [31:0] btbMeta_9; // @[bht.scala 114:26]
  reg [31:0] btbMeta_10; // @[bht.scala 114:26]
  reg [31:0] btbMeta_11; // @[bht.scala 114:26]
  reg [31:0] btbMeta_12; // @[bht.scala 114:26]
  reg [31:0] btbMeta_13; // @[bht.scala 114:26]
  reg [31:0] btbMeta_14; // @[bht.scala 114:26]
  reg [31:0] btbMeta_15; // @[bht.scala 114:26]
  reg [31:0] btbMeta_16; // @[bht.scala 114:26]
  reg [31:0] btbMeta_17; // @[bht.scala 114:26]
  reg [31:0] btbMeta_18; // @[bht.scala 114:26]
  reg [31:0] btbMeta_19; // @[bht.scala 114:26]
  reg [31:0] btbMeta_20; // @[bht.scala 114:26]
  reg [31:0] btbMeta_21; // @[bht.scala 114:26]
  reg [31:0] btbMeta_22; // @[bht.scala 114:26]
  reg [31:0] btbMeta_23; // @[bht.scala 114:26]
  reg [31:0] btbMeta_24; // @[bht.scala 114:26]
  reg [31:0] btbMeta_25; // @[bht.scala 114:26]
  reg [31:0] btbMeta_26; // @[bht.scala 114:26]
  reg [31:0] btbMeta_27; // @[bht.scala 114:26]
  reg [31:0] btbMeta_28; // @[bht.scala 114:26]
  reg [31:0] btbMeta_29; // @[bht.scala 114:26]
  reg [31:0] btbMeta_30; // @[bht.scala 114:26]
  reg [31:0] btbMeta_31; // @[bht.scala 114:26]
  reg [31:0] btbMeta_32; // @[bht.scala 114:26]
  reg [31:0] btbMeta_33; // @[bht.scala 114:26]
  reg [31:0] btbMeta_34; // @[bht.scala 114:26]
  reg [31:0] btbMeta_35; // @[bht.scala 114:26]
  reg [31:0] btbMeta_36; // @[bht.scala 114:26]
  reg [31:0] btbMeta_37; // @[bht.scala 114:26]
  reg [31:0] btbMeta_38; // @[bht.scala 114:26]
  reg [31:0] btbMeta_39; // @[bht.scala 114:26]
  reg [31:0] btbMeta_40; // @[bht.scala 114:26]
  reg [31:0] btbMeta_41; // @[bht.scala 114:26]
  reg [31:0] btbMeta_42; // @[bht.scala 114:26]
  reg [31:0] btbMeta_43; // @[bht.scala 114:26]
  reg [31:0] btbMeta_44; // @[bht.scala 114:26]
  reg [31:0] btbMeta_45; // @[bht.scala 114:26]
  reg [31:0] btbMeta_46; // @[bht.scala 114:26]
  reg [31:0] btbMeta_47; // @[bht.scala 114:26]
  reg [31:0] btbMeta_48; // @[bht.scala 114:26]
  reg [31:0] btbMeta_49; // @[bht.scala 114:26]
  reg [31:0] btbMeta_50; // @[bht.scala 114:26]
  reg [31:0] btbMeta_51; // @[bht.scala 114:26]
  reg [31:0] btbMeta_52; // @[bht.scala 114:26]
  reg [31:0] btbMeta_53; // @[bht.scala 114:26]
  reg [31:0] btbMeta_54; // @[bht.scala 114:26]
  reg [31:0] btbMeta_55; // @[bht.scala 114:26]
  reg [31:0] btbMeta_56; // @[bht.scala 114:26]
  reg [31:0] btbMeta_57; // @[bht.scala 114:26]
  reg [31:0] btbMeta_58; // @[bht.scala 114:26]
  reg [31:0] btbMeta_59; // @[bht.scala 114:26]
  reg [31:0] btbMeta_60; // @[bht.scala 114:26]
  reg [31:0] btbMeta_61; // @[bht.scala 114:26]
  reg [31:0] btbMeta_62; // @[bht.scala 114:26]
  reg [31:0] btbMeta_63; // @[bht.scala 114:26]
  reg [31:0] btbMeta_64; // @[bht.scala 114:26]
  reg [31:0] btbMeta_65; // @[bht.scala 114:26]
  reg [31:0] btbMeta_66; // @[bht.scala 114:26]
  reg [31:0] btbMeta_67; // @[bht.scala 114:26]
  reg [31:0] btbMeta_68; // @[bht.scala 114:26]
  reg [31:0] btbMeta_69; // @[bht.scala 114:26]
  reg [31:0] btbMeta_70; // @[bht.scala 114:26]
  reg [31:0] btbMeta_71; // @[bht.scala 114:26]
  reg [31:0] btbMeta_72; // @[bht.scala 114:26]
  reg [31:0] btbMeta_73; // @[bht.scala 114:26]
  reg [31:0] btbMeta_74; // @[bht.scala 114:26]
  reg [31:0] btbMeta_75; // @[bht.scala 114:26]
  reg [31:0] btbMeta_76; // @[bht.scala 114:26]
  reg [31:0] btbMeta_77; // @[bht.scala 114:26]
  reg [31:0] btbMeta_78; // @[bht.scala 114:26]
  reg [31:0] btbMeta_79; // @[bht.scala 114:26]
  reg [31:0] btbMeta_80; // @[bht.scala 114:26]
  reg [31:0] btbMeta_81; // @[bht.scala 114:26]
  reg [31:0] btbMeta_82; // @[bht.scala 114:26]
  reg [31:0] btbMeta_83; // @[bht.scala 114:26]
  reg [31:0] btbMeta_84; // @[bht.scala 114:26]
  reg [31:0] btbMeta_85; // @[bht.scala 114:26]
  reg [31:0] btbMeta_86; // @[bht.scala 114:26]
  reg [31:0] btbMeta_87; // @[bht.scala 114:26]
  reg [31:0] btbMeta_88; // @[bht.scala 114:26]
  reg [31:0] btbMeta_89; // @[bht.scala 114:26]
  reg [31:0] btbMeta_90; // @[bht.scala 114:26]
  reg [31:0] btbMeta_91; // @[bht.scala 114:26]
  reg [31:0] btbMeta_92; // @[bht.scala 114:26]
  reg [31:0] btbMeta_93; // @[bht.scala 114:26]
  reg [31:0] btbMeta_94; // @[bht.scala 114:26]
  reg [31:0] btbMeta_95; // @[bht.scala 114:26]
  reg [31:0] btbMeta_96; // @[bht.scala 114:26]
  reg [31:0] btbMeta_97; // @[bht.scala 114:26]
  reg [31:0] btbMeta_98; // @[bht.scala 114:26]
  reg [31:0] btbMeta_99; // @[bht.scala 114:26]
  reg [31:0] btbMeta_100; // @[bht.scala 114:26]
  reg [31:0] btbMeta_101; // @[bht.scala 114:26]
  reg [31:0] btbMeta_102; // @[bht.scala 114:26]
  reg [31:0] btbMeta_103; // @[bht.scala 114:26]
  reg [31:0] btbMeta_104; // @[bht.scala 114:26]
  reg [31:0] btbMeta_105; // @[bht.scala 114:26]
  reg [31:0] btbMeta_106; // @[bht.scala 114:26]
  reg [31:0] btbMeta_107; // @[bht.scala 114:26]
  reg [31:0] btbMeta_108; // @[bht.scala 114:26]
  reg [31:0] btbMeta_109; // @[bht.scala 114:26]
  reg [31:0] btbMeta_110; // @[bht.scala 114:26]
  reg [31:0] btbMeta_111; // @[bht.scala 114:26]
  reg [31:0] btbMeta_112; // @[bht.scala 114:26]
  reg [31:0] btbMeta_113; // @[bht.scala 114:26]
  reg [31:0] btbMeta_114; // @[bht.scala 114:26]
  reg [31:0] btbMeta_115; // @[bht.scala 114:26]
  reg [31:0] btbMeta_116; // @[bht.scala 114:26]
  reg [31:0] btbMeta_117; // @[bht.scala 114:26]
  reg [31:0] btbMeta_118; // @[bht.scala 114:26]
  reg [31:0] btbMeta_119; // @[bht.scala 114:26]
  reg [31:0] btbMeta_120; // @[bht.scala 114:26]
  reg [31:0] btbMeta_121; // @[bht.scala 114:26]
  reg [31:0] btbMeta_122; // @[bht.scala 114:26]
  reg [31:0] btbMeta_123; // @[bht.scala 114:26]
  reg [31:0] btbMeta_124; // @[bht.scala 114:26]
  reg [31:0] btbMeta_125; // @[bht.scala 114:26]
  reg [31:0] btbMeta_126; // @[bht.scala 114:26]
  reg [31:0] btbMeta_127; // @[bht.scala 114:26]
  wire  p1Addr_hash0 = io_pc[2] ^ io_pc[14]; // @[bht.scala 90:27]
  wire  _p1Addr_hash1_T_2 = io_pc[9] ^ io_pc[10]; // @[bht.scala 91:28]
  wire  p1Addr_hash1 = io_pc[9] ^ io_pc[10] ^ (io_pc[3] ^ io_pc[15]); // @[bht.scala 91:39]
  wire  p1Addr_hash2 = io_pc[4] ^ (io_pc[10] ^ io_pc[11]); // @[bht.scala 92:27]
  wire  p1Addr_hash3 = io_pc[5] ^ (io_pc[11] ^ io_pc[12]); // @[bht.scala 93:27]
  wire  p1Addr_hash4 = io_pc[6] ^ (io_pc[12] ^ io_pc[13]); // @[bht.scala 94:27]
  wire  p1Addr_hash5 = io_pc[7] ^ (io_pc[13] ^ io_pc[14]); // @[bht.scala 95:27]
  wire  p1Addr_hash6 = io_pc[8] ^ _p1Addr_hash1_T_2; // @[bht.scala 96:27]
  wire [6:0] _p1Addr_T_6 = {p1Addr_hash6,p1Addr_hash5,p1Addr_hash4,p1Addr_hash3,p1Addr_hash2,p1Addr_hash1,p1Addr_hash0}; // @[bht.scala 97:58]
  wire [6:0] p1Addr = _p1Addr_T_6 ^ ghr; // @[bht.scala 102:26]
  wire [6:0] _GEN_1 = 7'h1 == _p1Addr_T_6 ? bht_1 : bht_0; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_2 = 7'h2 == _p1Addr_T_6 ? bht_2 : _GEN_1; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_3 = 7'h3 == _p1Addr_T_6 ? bht_3 : _GEN_2; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_4 = 7'h4 == _p1Addr_T_6 ? bht_4 : _GEN_3; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_5 = 7'h5 == _p1Addr_T_6 ? bht_5 : _GEN_4; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_6 = 7'h6 == _p1Addr_T_6 ? bht_6 : _GEN_5; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_7 = 7'h7 == _p1Addr_T_6 ? bht_7 : _GEN_6; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_8 = 7'h8 == _p1Addr_T_6 ? bht_8 : _GEN_7; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_9 = 7'h9 == _p1Addr_T_6 ? bht_9 : _GEN_8; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_10 = 7'ha == _p1Addr_T_6 ? bht_10 : _GEN_9; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_11 = 7'hb == _p1Addr_T_6 ? bht_11 : _GEN_10; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_12 = 7'hc == _p1Addr_T_6 ? bht_12 : _GEN_11; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_13 = 7'hd == _p1Addr_T_6 ? bht_13 : _GEN_12; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_14 = 7'he == _p1Addr_T_6 ? bht_14 : _GEN_13; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_15 = 7'hf == _p1Addr_T_6 ? bht_15 : _GEN_14; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_16 = 7'h10 == _p1Addr_T_6 ? bht_16 : _GEN_15; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_17 = 7'h11 == _p1Addr_T_6 ? bht_17 : _GEN_16; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_18 = 7'h12 == _p1Addr_T_6 ? bht_18 : _GEN_17; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_19 = 7'h13 == _p1Addr_T_6 ? bht_19 : _GEN_18; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_20 = 7'h14 == _p1Addr_T_6 ? bht_20 : _GEN_19; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_21 = 7'h15 == _p1Addr_T_6 ? bht_21 : _GEN_20; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_22 = 7'h16 == _p1Addr_T_6 ? bht_22 : _GEN_21; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_23 = 7'h17 == _p1Addr_T_6 ? bht_23 : _GEN_22; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_24 = 7'h18 == _p1Addr_T_6 ? bht_24 : _GEN_23; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_25 = 7'h19 == _p1Addr_T_6 ? bht_25 : _GEN_24; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_26 = 7'h1a == _p1Addr_T_6 ? bht_26 : _GEN_25; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_27 = 7'h1b == _p1Addr_T_6 ? bht_27 : _GEN_26; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_28 = 7'h1c == _p1Addr_T_6 ? bht_28 : _GEN_27; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_29 = 7'h1d == _p1Addr_T_6 ? bht_29 : _GEN_28; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_30 = 7'h1e == _p1Addr_T_6 ? bht_30 : _GEN_29; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_31 = 7'h1f == _p1Addr_T_6 ? bht_31 : _GEN_30; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_32 = 7'h20 == _p1Addr_T_6 ? bht_32 : _GEN_31; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_33 = 7'h21 == _p1Addr_T_6 ? bht_33 : _GEN_32; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_34 = 7'h22 == _p1Addr_T_6 ? bht_34 : _GEN_33; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_35 = 7'h23 == _p1Addr_T_6 ? bht_35 : _GEN_34; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_36 = 7'h24 == _p1Addr_T_6 ? bht_36 : _GEN_35; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_37 = 7'h25 == _p1Addr_T_6 ? bht_37 : _GEN_36; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_38 = 7'h26 == _p1Addr_T_6 ? bht_38 : _GEN_37; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_39 = 7'h27 == _p1Addr_T_6 ? bht_39 : _GEN_38; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_40 = 7'h28 == _p1Addr_T_6 ? bht_40 : _GEN_39; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_41 = 7'h29 == _p1Addr_T_6 ? bht_41 : _GEN_40; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_42 = 7'h2a == _p1Addr_T_6 ? bht_42 : _GEN_41; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_43 = 7'h2b == _p1Addr_T_6 ? bht_43 : _GEN_42; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_44 = 7'h2c == _p1Addr_T_6 ? bht_44 : _GEN_43; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_45 = 7'h2d == _p1Addr_T_6 ? bht_45 : _GEN_44; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_46 = 7'h2e == _p1Addr_T_6 ? bht_46 : _GEN_45; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_47 = 7'h2f == _p1Addr_T_6 ? bht_47 : _GEN_46; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_48 = 7'h30 == _p1Addr_T_6 ? bht_48 : _GEN_47; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_49 = 7'h31 == _p1Addr_T_6 ? bht_49 : _GEN_48; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_50 = 7'h32 == _p1Addr_T_6 ? bht_50 : _GEN_49; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_51 = 7'h33 == _p1Addr_T_6 ? bht_51 : _GEN_50; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_52 = 7'h34 == _p1Addr_T_6 ? bht_52 : _GEN_51; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_53 = 7'h35 == _p1Addr_T_6 ? bht_53 : _GEN_52; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_54 = 7'h36 == _p1Addr_T_6 ? bht_54 : _GEN_53; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_55 = 7'h37 == _p1Addr_T_6 ? bht_55 : _GEN_54; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_56 = 7'h38 == _p1Addr_T_6 ? bht_56 : _GEN_55; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_57 = 7'h39 == _p1Addr_T_6 ? bht_57 : _GEN_56; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_58 = 7'h3a == _p1Addr_T_6 ? bht_58 : _GEN_57; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_59 = 7'h3b == _p1Addr_T_6 ? bht_59 : _GEN_58; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_60 = 7'h3c == _p1Addr_T_6 ? bht_60 : _GEN_59; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_61 = 7'h3d == _p1Addr_T_6 ? bht_61 : _GEN_60; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_62 = 7'h3e == _p1Addr_T_6 ? bht_62 : _GEN_61; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_63 = 7'h3f == _p1Addr_T_6 ? bht_63 : _GEN_62; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_64 = 7'h40 == _p1Addr_T_6 ? bht_64 : _GEN_63; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_65 = 7'h41 == _p1Addr_T_6 ? bht_65 : _GEN_64; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_66 = 7'h42 == _p1Addr_T_6 ? bht_66 : _GEN_65; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_67 = 7'h43 == _p1Addr_T_6 ? bht_67 : _GEN_66; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_68 = 7'h44 == _p1Addr_T_6 ? bht_68 : _GEN_67; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_69 = 7'h45 == _p1Addr_T_6 ? bht_69 : _GEN_68; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_70 = 7'h46 == _p1Addr_T_6 ? bht_70 : _GEN_69; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_71 = 7'h47 == _p1Addr_T_6 ? bht_71 : _GEN_70; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_72 = 7'h48 == _p1Addr_T_6 ? bht_72 : _GEN_71; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_73 = 7'h49 == _p1Addr_T_6 ? bht_73 : _GEN_72; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_74 = 7'h4a == _p1Addr_T_6 ? bht_74 : _GEN_73; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_75 = 7'h4b == _p1Addr_T_6 ? bht_75 : _GEN_74; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_76 = 7'h4c == _p1Addr_T_6 ? bht_76 : _GEN_75; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_77 = 7'h4d == _p1Addr_T_6 ? bht_77 : _GEN_76; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_78 = 7'h4e == _p1Addr_T_6 ? bht_78 : _GEN_77; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_79 = 7'h4f == _p1Addr_T_6 ? bht_79 : _GEN_78; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_80 = 7'h50 == _p1Addr_T_6 ? bht_80 : _GEN_79; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_81 = 7'h51 == _p1Addr_T_6 ? bht_81 : _GEN_80; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_82 = 7'h52 == _p1Addr_T_6 ? bht_82 : _GEN_81; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_83 = 7'h53 == _p1Addr_T_6 ? bht_83 : _GEN_82; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_84 = 7'h54 == _p1Addr_T_6 ? bht_84 : _GEN_83; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_85 = 7'h55 == _p1Addr_T_6 ? bht_85 : _GEN_84; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_86 = 7'h56 == _p1Addr_T_6 ? bht_86 : _GEN_85; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_87 = 7'h57 == _p1Addr_T_6 ? bht_87 : _GEN_86; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_88 = 7'h58 == _p1Addr_T_6 ? bht_88 : _GEN_87; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_89 = 7'h59 == _p1Addr_T_6 ? bht_89 : _GEN_88; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_90 = 7'h5a == _p1Addr_T_6 ? bht_90 : _GEN_89; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_91 = 7'h5b == _p1Addr_T_6 ? bht_91 : _GEN_90; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_92 = 7'h5c == _p1Addr_T_6 ? bht_92 : _GEN_91; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_93 = 7'h5d == _p1Addr_T_6 ? bht_93 : _GEN_92; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_94 = 7'h5e == _p1Addr_T_6 ? bht_94 : _GEN_93; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_95 = 7'h5f == _p1Addr_T_6 ? bht_95 : _GEN_94; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_96 = 7'h60 == _p1Addr_T_6 ? bht_96 : _GEN_95; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_97 = 7'h61 == _p1Addr_T_6 ? bht_97 : _GEN_96; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_98 = 7'h62 == _p1Addr_T_6 ? bht_98 : _GEN_97; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_99 = 7'h63 == _p1Addr_T_6 ? bht_99 : _GEN_98; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_100 = 7'h64 == _p1Addr_T_6 ? bht_100 : _GEN_99; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_101 = 7'h65 == _p1Addr_T_6 ? bht_101 : _GEN_100; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_102 = 7'h66 == _p1Addr_T_6 ? bht_102 : _GEN_101; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_103 = 7'h67 == _p1Addr_T_6 ? bht_103 : _GEN_102; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_104 = 7'h68 == _p1Addr_T_6 ? bht_104 : _GEN_103; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_105 = 7'h69 == _p1Addr_T_6 ? bht_105 : _GEN_104; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_106 = 7'h6a == _p1Addr_T_6 ? bht_106 : _GEN_105; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_107 = 7'h6b == _p1Addr_T_6 ? bht_107 : _GEN_106; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_108 = 7'h6c == _p1Addr_T_6 ? bht_108 : _GEN_107; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_109 = 7'h6d == _p1Addr_T_6 ? bht_109 : _GEN_108; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_110 = 7'h6e == _p1Addr_T_6 ? bht_110 : _GEN_109; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_111 = 7'h6f == _p1Addr_T_6 ? bht_111 : _GEN_110; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_112 = 7'h70 == _p1Addr_T_6 ? bht_112 : _GEN_111; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_113 = 7'h71 == _p1Addr_T_6 ? bht_113 : _GEN_112; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_114 = 7'h72 == _p1Addr_T_6 ? bht_114 : _GEN_113; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_115 = 7'h73 == _p1Addr_T_6 ? bht_115 : _GEN_114; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_116 = 7'h74 == _p1Addr_T_6 ? bht_116 : _GEN_115; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_117 = 7'h75 == _p1Addr_T_6 ? bht_117 : _GEN_116; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_118 = 7'h76 == _p1Addr_T_6 ? bht_118 : _GEN_117; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_119 = 7'h77 == _p1Addr_T_6 ? bht_119 : _GEN_118; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_120 = 7'h78 == _p1Addr_T_6 ? bht_120 : _GEN_119; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_121 = 7'h79 == _p1Addr_T_6 ? bht_121 : _GEN_120; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_122 = 7'h7a == _p1Addr_T_6 ? bht_122 : _GEN_121; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_123 = 7'h7b == _p1Addr_T_6 ? bht_123 : _GEN_122; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_124 = 7'h7c == _p1Addr_T_6 ? bht_124 : _GEN_123; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_125 = 7'h7d == _p1Addr_T_6 ? bht_125 : _GEN_124; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_126 = 7'h7e == _p1Addr_T_6 ? bht_126 : _GEN_125; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_127 = 7'h7f == _p1Addr_T_6 ? bht_127 : _GEN_126; // @[bht.scala 102:{26,26}]
  wire [6:0] _pht2Data_T_7 = _p1Addr_T_6 ^ _GEN_127; // @[bht.scala 102:26]
  wire [1:0] _GEN_129 = 7'h1 == p1Addr ? pht_0_1 : pht_0_0; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_130 = 7'h2 == p1Addr ? pht_0_2 : _GEN_129; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_131 = 7'h3 == p1Addr ? pht_0_3 : _GEN_130; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_132 = 7'h4 == p1Addr ? pht_0_4 : _GEN_131; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_133 = 7'h5 == p1Addr ? pht_0_5 : _GEN_132; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_134 = 7'h6 == p1Addr ? pht_0_6 : _GEN_133; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_135 = 7'h7 == p1Addr ? pht_0_7 : _GEN_134; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_136 = 7'h8 == p1Addr ? pht_0_8 : _GEN_135; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_137 = 7'h9 == p1Addr ? pht_0_9 : _GEN_136; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_138 = 7'ha == p1Addr ? pht_0_10 : _GEN_137; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_139 = 7'hb == p1Addr ? pht_0_11 : _GEN_138; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_140 = 7'hc == p1Addr ? pht_0_12 : _GEN_139; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_141 = 7'hd == p1Addr ? pht_0_13 : _GEN_140; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_142 = 7'he == p1Addr ? pht_0_14 : _GEN_141; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_143 = 7'hf == p1Addr ? pht_0_15 : _GEN_142; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_144 = 7'h10 == p1Addr ? pht_0_16 : _GEN_143; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_145 = 7'h11 == p1Addr ? pht_0_17 : _GEN_144; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_146 = 7'h12 == p1Addr ? pht_0_18 : _GEN_145; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_147 = 7'h13 == p1Addr ? pht_0_19 : _GEN_146; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_148 = 7'h14 == p1Addr ? pht_0_20 : _GEN_147; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_149 = 7'h15 == p1Addr ? pht_0_21 : _GEN_148; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_150 = 7'h16 == p1Addr ? pht_0_22 : _GEN_149; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_151 = 7'h17 == p1Addr ? pht_0_23 : _GEN_150; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_152 = 7'h18 == p1Addr ? pht_0_24 : _GEN_151; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_153 = 7'h19 == p1Addr ? pht_0_25 : _GEN_152; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_154 = 7'h1a == p1Addr ? pht_0_26 : _GEN_153; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_155 = 7'h1b == p1Addr ? pht_0_27 : _GEN_154; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_156 = 7'h1c == p1Addr ? pht_0_28 : _GEN_155; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_157 = 7'h1d == p1Addr ? pht_0_29 : _GEN_156; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_158 = 7'h1e == p1Addr ? pht_0_30 : _GEN_157; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_159 = 7'h1f == p1Addr ? pht_0_31 : _GEN_158; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_160 = 7'h20 == p1Addr ? pht_0_32 : _GEN_159; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_161 = 7'h21 == p1Addr ? pht_0_33 : _GEN_160; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_162 = 7'h22 == p1Addr ? pht_0_34 : _GEN_161; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_163 = 7'h23 == p1Addr ? pht_0_35 : _GEN_162; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_164 = 7'h24 == p1Addr ? pht_0_36 : _GEN_163; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_165 = 7'h25 == p1Addr ? pht_0_37 : _GEN_164; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_166 = 7'h26 == p1Addr ? pht_0_38 : _GEN_165; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_167 = 7'h27 == p1Addr ? pht_0_39 : _GEN_166; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_168 = 7'h28 == p1Addr ? pht_0_40 : _GEN_167; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_169 = 7'h29 == p1Addr ? pht_0_41 : _GEN_168; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_170 = 7'h2a == p1Addr ? pht_0_42 : _GEN_169; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_171 = 7'h2b == p1Addr ? pht_0_43 : _GEN_170; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_172 = 7'h2c == p1Addr ? pht_0_44 : _GEN_171; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_173 = 7'h2d == p1Addr ? pht_0_45 : _GEN_172; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_174 = 7'h2e == p1Addr ? pht_0_46 : _GEN_173; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_175 = 7'h2f == p1Addr ? pht_0_47 : _GEN_174; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_176 = 7'h30 == p1Addr ? pht_0_48 : _GEN_175; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_177 = 7'h31 == p1Addr ? pht_0_49 : _GEN_176; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_178 = 7'h32 == p1Addr ? pht_0_50 : _GEN_177; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_179 = 7'h33 == p1Addr ? pht_0_51 : _GEN_178; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_180 = 7'h34 == p1Addr ? pht_0_52 : _GEN_179; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_181 = 7'h35 == p1Addr ? pht_0_53 : _GEN_180; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_182 = 7'h36 == p1Addr ? pht_0_54 : _GEN_181; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_183 = 7'h37 == p1Addr ? pht_0_55 : _GEN_182; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_184 = 7'h38 == p1Addr ? pht_0_56 : _GEN_183; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_185 = 7'h39 == p1Addr ? pht_0_57 : _GEN_184; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_186 = 7'h3a == p1Addr ? pht_0_58 : _GEN_185; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_187 = 7'h3b == p1Addr ? pht_0_59 : _GEN_186; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_188 = 7'h3c == p1Addr ? pht_0_60 : _GEN_187; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_189 = 7'h3d == p1Addr ? pht_0_61 : _GEN_188; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_190 = 7'h3e == p1Addr ? pht_0_62 : _GEN_189; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_191 = 7'h3f == p1Addr ? pht_0_63 : _GEN_190; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_192 = 7'h40 == p1Addr ? pht_0_64 : _GEN_191; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_193 = 7'h41 == p1Addr ? pht_0_65 : _GEN_192; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_194 = 7'h42 == p1Addr ? pht_0_66 : _GEN_193; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_195 = 7'h43 == p1Addr ? pht_0_67 : _GEN_194; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_196 = 7'h44 == p1Addr ? pht_0_68 : _GEN_195; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_197 = 7'h45 == p1Addr ? pht_0_69 : _GEN_196; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_198 = 7'h46 == p1Addr ? pht_0_70 : _GEN_197; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_199 = 7'h47 == p1Addr ? pht_0_71 : _GEN_198; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_200 = 7'h48 == p1Addr ? pht_0_72 : _GEN_199; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_201 = 7'h49 == p1Addr ? pht_0_73 : _GEN_200; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_202 = 7'h4a == p1Addr ? pht_0_74 : _GEN_201; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_203 = 7'h4b == p1Addr ? pht_0_75 : _GEN_202; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_204 = 7'h4c == p1Addr ? pht_0_76 : _GEN_203; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_205 = 7'h4d == p1Addr ? pht_0_77 : _GEN_204; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_206 = 7'h4e == p1Addr ? pht_0_78 : _GEN_205; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_207 = 7'h4f == p1Addr ? pht_0_79 : _GEN_206; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_208 = 7'h50 == p1Addr ? pht_0_80 : _GEN_207; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_209 = 7'h51 == p1Addr ? pht_0_81 : _GEN_208; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_210 = 7'h52 == p1Addr ? pht_0_82 : _GEN_209; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_211 = 7'h53 == p1Addr ? pht_0_83 : _GEN_210; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_212 = 7'h54 == p1Addr ? pht_0_84 : _GEN_211; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_213 = 7'h55 == p1Addr ? pht_0_85 : _GEN_212; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_214 = 7'h56 == p1Addr ? pht_0_86 : _GEN_213; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_215 = 7'h57 == p1Addr ? pht_0_87 : _GEN_214; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_216 = 7'h58 == p1Addr ? pht_0_88 : _GEN_215; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_217 = 7'h59 == p1Addr ? pht_0_89 : _GEN_216; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_218 = 7'h5a == p1Addr ? pht_0_90 : _GEN_217; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_219 = 7'h5b == p1Addr ? pht_0_91 : _GEN_218; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_220 = 7'h5c == p1Addr ? pht_0_92 : _GEN_219; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_221 = 7'h5d == p1Addr ? pht_0_93 : _GEN_220; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_222 = 7'h5e == p1Addr ? pht_0_94 : _GEN_221; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_223 = 7'h5f == p1Addr ? pht_0_95 : _GEN_222; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_224 = 7'h60 == p1Addr ? pht_0_96 : _GEN_223; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_225 = 7'h61 == p1Addr ? pht_0_97 : _GEN_224; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_226 = 7'h62 == p1Addr ? pht_0_98 : _GEN_225; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_227 = 7'h63 == p1Addr ? pht_0_99 : _GEN_226; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_228 = 7'h64 == p1Addr ? pht_0_100 : _GEN_227; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_229 = 7'h65 == p1Addr ? pht_0_101 : _GEN_228; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_230 = 7'h66 == p1Addr ? pht_0_102 : _GEN_229; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_231 = 7'h67 == p1Addr ? pht_0_103 : _GEN_230; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_232 = 7'h68 == p1Addr ? pht_0_104 : _GEN_231; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_233 = 7'h69 == p1Addr ? pht_0_105 : _GEN_232; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_234 = 7'h6a == p1Addr ? pht_0_106 : _GEN_233; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_235 = 7'h6b == p1Addr ? pht_0_107 : _GEN_234; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_236 = 7'h6c == p1Addr ? pht_0_108 : _GEN_235; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_237 = 7'h6d == p1Addr ? pht_0_109 : _GEN_236; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_238 = 7'h6e == p1Addr ? pht_0_110 : _GEN_237; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_239 = 7'h6f == p1Addr ? pht_0_111 : _GEN_238; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_240 = 7'h70 == p1Addr ? pht_0_112 : _GEN_239; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_241 = 7'h71 == p1Addr ? pht_0_113 : _GEN_240; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_242 = 7'h72 == p1Addr ? pht_0_114 : _GEN_241; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_243 = 7'h73 == p1Addr ? pht_0_115 : _GEN_242; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_244 = 7'h74 == p1Addr ? pht_0_116 : _GEN_243; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_245 = 7'h75 == p1Addr ? pht_0_117 : _GEN_244; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_246 = 7'h76 == p1Addr ? pht_0_118 : _GEN_245; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_247 = 7'h77 == p1Addr ? pht_0_119 : _GEN_246; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_248 = 7'h78 == p1Addr ? pht_0_120 : _GEN_247; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_249 = 7'h79 == p1Addr ? pht_0_121 : _GEN_248; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_250 = 7'h7a == p1Addr ? pht_0_122 : _GEN_249; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_251 = 7'h7b == p1Addr ? pht_0_123 : _GEN_250; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_252 = 7'h7c == p1Addr ? pht_0_124 : _GEN_251; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_253 = 7'h7d == p1Addr ? pht_0_125 : _GEN_252; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_254 = 7'h7e == p1Addr ? pht_0_126 : _GEN_253; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_255 = 7'h7f == p1Addr ? pht_0_127 : _GEN_254; // @[bht.scala 123:{32,32}]
  wire [1:0] _GEN_257 = 7'h1 == _pht2Data_T_7 ? pht_2_1 : pht_2_0; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_258 = 7'h2 == _pht2Data_T_7 ? pht_2_2 : _GEN_257; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_259 = 7'h3 == _pht2Data_T_7 ? pht_2_3 : _GEN_258; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_260 = 7'h4 == _pht2Data_T_7 ? pht_2_4 : _GEN_259; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_261 = 7'h5 == _pht2Data_T_7 ? pht_2_5 : _GEN_260; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_262 = 7'h6 == _pht2Data_T_7 ? pht_2_6 : _GEN_261; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_263 = 7'h7 == _pht2Data_T_7 ? pht_2_7 : _GEN_262; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_264 = 7'h8 == _pht2Data_T_7 ? pht_2_8 : _GEN_263; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_265 = 7'h9 == _pht2Data_T_7 ? pht_2_9 : _GEN_264; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_266 = 7'ha == _pht2Data_T_7 ? pht_2_10 : _GEN_265; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_267 = 7'hb == _pht2Data_T_7 ? pht_2_11 : _GEN_266; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_268 = 7'hc == _pht2Data_T_7 ? pht_2_12 : _GEN_267; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_269 = 7'hd == _pht2Data_T_7 ? pht_2_13 : _GEN_268; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_270 = 7'he == _pht2Data_T_7 ? pht_2_14 : _GEN_269; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_271 = 7'hf == _pht2Data_T_7 ? pht_2_15 : _GEN_270; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_272 = 7'h10 == _pht2Data_T_7 ? pht_2_16 : _GEN_271; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_273 = 7'h11 == _pht2Data_T_7 ? pht_2_17 : _GEN_272; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_274 = 7'h12 == _pht2Data_T_7 ? pht_2_18 : _GEN_273; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_275 = 7'h13 == _pht2Data_T_7 ? pht_2_19 : _GEN_274; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_276 = 7'h14 == _pht2Data_T_7 ? pht_2_20 : _GEN_275; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_277 = 7'h15 == _pht2Data_T_7 ? pht_2_21 : _GEN_276; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_278 = 7'h16 == _pht2Data_T_7 ? pht_2_22 : _GEN_277; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_279 = 7'h17 == _pht2Data_T_7 ? pht_2_23 : _GEN_278; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_280 = 7'h18 == _pht2Data_T_7 ? pht_2_24 : _GEN_279; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_281 = 7'h19 == _pht2Data_T_7 ? pht_2_25 : _GEN_280; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_282 = 7'h1a == _pht2Data_T_7 ? pht_2_26 : _GEN_281; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_283 = 7'h1b == _pht2Data_T_7 ? pht_2_27 : _GEN_282; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_284 = 7'h1c == _pht2Data_T_7 ? pht_2_28 : _GEN_283; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_285 = 7'h1d == _pht2Data_T_7 ? pht_2_29 : _GEN_284; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_286 = 7'h1e == _pht2Data_T_7 ? pht_2_30 : _GEN_285; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_287 = 7'h1f == _pht2Data_T_7 ? pht_2_31 : _GEN_286; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_288 = 7'h20 == _pht2Data_T_7 ? pht_2_32 : _GEN_287; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_289 = 7'h21 == _pht2Data_T_7 ? pht_2_33 : _GEN_288; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_290 = 7'h22 == _pht2Data_T_7 ? pht_2_34 : _GEN_289; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_291 = 7'h23 == _pht2Data_T_7 ? pht_2_35 : _GEN_290; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_292 = 7'h24 == _pht2Data_T_7 ? pht_2_36 : _GEN_291; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_293 = 7'h25 == _pht2Data_T_7 ? pht_2_37 : _GEN_292; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_294 = 7'h26 == _pht2Data_T_7 ? pht_2_38 : _GEN_293; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_295 = 7'h27 == _pht2Data_T_7 ? pht_2_39 : _GEN_294; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_296 = 7'h28 == _pht2Data_T_7 ? pht_2_40 : _GEN_295; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_297 = 7'h29 == _pht2Data_T_7 ? pht_2_41 : _GEN_296; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_298 = 7'h2a == _pht2Data_T_7 ? pht_2_42 : _GEN_297; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_299 = 7'h2b == _pht2Data_T_7 ? pht_2_43 : _GEN_298; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_300 = 7'h2c == _pht2Data_T_7 ? pht_2_44 : _GEN_299; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_301 = 7'h2d == _pht2Data_T_7 ? pht_2_45 : _GEN_300; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_302 = 7'h2e == _pht2Data_T_7 ? pht_2_46 : _GEN_301; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_303 = 7'h2f == _pht2Data_T_7 ? pht_2_47 : _GEN_302; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_304 = 7'h30 == _pht2Data_T_7 ? pht_2_48 : _GEN_303; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_305 = 7'h31 == _pht2Data_T_7 ? pht_2_49 : _GEN_304; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_306 = 7'h32 == _pht2Data_T_7 ? pht_2_50 : _GEN_305; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_307 = 7'h33 == _pht2Data_T_7 ? pht_2_51 : _GEN_306; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_308 = 7'h34 == _pht2Data_T_7 ? pht_2_52 : _GEN_307; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_309 = 7'h35 == _pht2Data_T_7 ? pht_2_53 : _GEN_308; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_310 = 7'h36 == _pht2Data_T_7 ? pht_2_54 : _GEN_309; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_311 = 7'h37 == _pht2Data_T_7 ? pht_2_55 : _GEN_310; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_312 = 7'h38 == _pht2Data_T_7 ? pht_2_56 : _GEN_311; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_313 = 7'h39 == _pht2Data_T_7 ? pht_2_57 : _GEN_312; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_314 = 7'h3a == _pht2Data_T_7 ? pht_2_58 : _GEN_313; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_315 = 7'h3b == _pht2Data_T_7 ? pht_2_59 : _GEN_314; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_316 = 7'h3c == _pht2Data_T_7 ? pht_2_60 : _GEN_315; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_317 = 7'h3d == _pht2Data_T_7 ? pht_2_61 : _GEN_316; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_318 = 7'h3e == _pht2Data_T_7 ? pht_2_62 : _GEN_317; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_319 = 7'h3f == _pht2Data_T_7 ? pht_2_63 : _GEN_318; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_320 = 7'h40 == _pht2Data_T_7 ? pht_2_64 : _GEN_319; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_321 = 7'h41 == _pht2Data_T_7 ? pht_2_65 : _GEN_320; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_322 = 7'h42 == _pht2Data_T_7 ? pht_2_66 : _GEN_321; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_323 = 7'h43 == _pht2Data_T_7 ? pht_2_67 : _GEN_322; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_324 = 7'h44 == _pht2Data_T_7 ? pht_2_68 : _GEN_323; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_325 = 7'h45 == _pht2Data_T_7 ? pht_2_69 : _GEN_324; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_326 = 7'h46 == _pht2Data_T_7 ? pht_2_70 : _GEN_325; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_327 = 7'h47 == _pht2Data_T_7 ? pht_2_71 : _GEN_326; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_328 = 7'h48 == _pht2Data_T_7 ? pht_2_72 : _GEN_327; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_329 = 7'h49 == _pht2Data_T_7 ? pht_2_73 : _GEN_328; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_330 = 7'h4a == _pht2Data_T_7 ? pht_2_74 : _GEN_329; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_331 = 7'h4b == _pht2Data_T_7 ? pht_2_75 : _GEN_330; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_332 = 7'h4c == _pht2Data_T_7 ? pht_2_76 : _GEN_331; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_333 = 7'h4d == _pht2Data_T_7 ? pht_2_77 : _GEN_332; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_334 = 7'h4e == _pht2Data_T_7 ? pht_2_78 : _GEN_333; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_335 = 7'h4f == _pht2Data_T_7 ? pht_2_79 : _GEN_334; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_336 = 7'h50 == _pht2Data_T_7 ? pht_2_80 : _GEN_335; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_337 = 7'h51 == _pht2Data_T_7 ? pht_2_81 : _GEN_336; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_338 = 7'h52 == _pht2Data_T_7 ? pht_2_82 : _GEN_337; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_339 = 7'h53 == _pht2Data_T_7 ? pht_2_83 : _GEN_338; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_340 = 7'h54 == _pht2Data_T_7 ? pht_2_84 : _GEN_339; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_341 = 7'h55 == _pht2Data_T_7 ? pht_2_85 : _GEN_340; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_342 = 7'h56 == _pht2Data_T_7 ? pht_2_86 : _GEN_341; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_343 = 7'h57 == _pht2Data_T_7 ? pht_2_87 : _GEN_342; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_344 = 7'h58 == _pht2Data_T_7 ? pht_2_88 : _GEN_343; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_345 = 7'h59 == _pht2Data_T_7 ? pht_2_89 : _GEN_344; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_346 = 7'h5a == _pht2Data_T_7 ? pht_2_90 : _GEN_345; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_347 = 7'h5b == _pht2Data_T_7 ? pht_2_91 : _GEN_346; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_348 = 7'h5c == _pht2Data_T_7 ? pht_2_92 : _GEN_347; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_349 = 7'h5d == _pht2Data_T_7 ? pht_2_93 : _GEN_348; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_350 = 7'h5e == _pht2Data_T_7 ? pht_2_94 : _GEN_349; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_351 = 7'h5f == _pht2Data_T_7 ? pht_2_95 : _GEN_350; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_352 = 7'h60 == _pht2Data_T_7 ? pht_2_96 : _GEN_351; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_353 = 7'h61 == _pht2Data_T_7 ? pht_2_97 : _GEN_352; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_354 = 7'h62 == _pht2Data_T_7 ? pht_2_98 : _GEN_353; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_355 = 7'h63 == _pht2Data_T_7 ? pht_2_99 : _GEN_354; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_356 = 7'h64 == _pht2Data_T_7 ? pht_2_100 : _GEN_355; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_357 = 7'h65 == _pht2Data_T_7 ? pht_2_101 : _GEN_356; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_358 = 7'h66 == _pht2Data_T_7 ? pht_2_102 : _GEN_357; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_359 = 7'h67 == _pht2Data_T_7 ? pht_2_103 : _GEN_358; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_360 = 7'h68 == _pht2Data_T_7 ? pht_2_104 : _GEN_359; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_361 = 7'h69 == _pht2Data_T_7 ? pht_2_105 : _GEN_360; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_362 = 7'h6a == _pht2Data_T_7 ? pht_2_106 : _GEN_361; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_363 = 7'h6b == _pht2Data_T_7 ? pht_2_107 : _GEN_362; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_364 = 7'h6c == _pht2Data_T_7 ? pht_2_108 : _GEN_363; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_365 = 7'h6d == _pht2Data_T_7 ? pht_2_109 : _GEN_364; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_366 = 7'h6e == _pht2Data_T_7 ? pht_2_110 : _GEN_365; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_367 = 7'h6f == _pht2Data_T_7 ? pht_2_111 : _GEN_366; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_368 = 7'h70 == _pht2Data_T_7 ? pht_2_112 : _GEN_367; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_369 = 7'h71 == _pht2Data_T_7 ? pht_2_113 : _GEN_368; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_370 = 7'h72 == _pht2Data_T_7 ? pht_2_114 : _GEN_369; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_371 = 7'h73 == _pht2Data_T_7 ? pht_2_115 : _GEN_370; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_372 = 7'h74 == _pht2Data_T_7 ? pht_2_116 : _GEN_371; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_373 = 7'h75 == _pht2Data_T_7 ? pht_2_117 : _GEN_372; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_374 = 7'h76 == _pht2Data_T_7 ? pht_2_118 : _GEN_373; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_375 = 7'h77 == _pht2Data_T_7 ? pht_2_119 : _GEN_374; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_376 = 7'h78 == _pht2Data_T_7 ? pht_2_120 : _GEN_375; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_377 = 7'h79 == _pht2Data_T_7 ? pht_2_121 : _GEN_376; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_378 = 7'h7a == _pht2Data_T_7 ? pht_2_122 : _GEN_377; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_379 = 7'h7b == _pht2Data_T_7 ? pht_2_123 : _GEN_378; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_380 = 7'h7c == _pht2Data_T_7 ? pht_2_124 : _GEN_379; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_381 = 7'h7d == _pht2Data_T_7 ? pht_2_125 : _GEN_380; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_382 = 7'h7e == _pht2Data_T_7 ? pht_2_126 : _GEN_381; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_383 = 7'h7f == _pht2Data_T_7 ? pht_2_127 : _GEN_382; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_385 = 7'h1 == p1Addr ? pht_1_1 : pht_1_0; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_386 = 7'h2 == p1Addr ? pht_1_2 : _GEN_385; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_387 = 7'h3 == p1Addr ? pht_1_3 : _GEN_386; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_388 = 7'h4 == p1Addr ? pht_1_4 : _GEN_387; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_389 = 7'h5 == p1Addr ? pht_1_5 : _GEN_388; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_390 = 7'h6 == p1Addr ? pht_1_6 : _GEN_389; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_391 = 7'h7 == p1Addr ? pht_1_7 : _GEN_390; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_392 = 7'h8 == p1Addr ? pht_1_8 : _GEN_391; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_393 = 7'h9 == p1Addr ? pht_1_9 : _GEN_392; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_394 = 7'ha == p1Addr ? pht_1_10 : _GEN_393; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_395 = 7'hb == p1Addr ? pht_1_11 : _GEN_394; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_396 = 7'hc == p1Addr ? pht_1_12 : _GEN_395; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_397 = 7'hd == p1Addr ? pht_1_13 : _GEN_396; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_398 = 7'he == p1Addr ? pht_1_14 : _GEN_397; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_399 = 7'hf == p1Addr ? pht_1_15 : _GEN_398; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_400 = 7'h10 == p1Addr ? pht_1_16 : _GEN_399; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_401 = 7'h11 == p1Addr ? pht_1_17 : _GEN_400; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_402 = 7'h12 == p1Addr ? pht_1_18 : _GEN_401; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_403 = 7'h13 == p1Addr ? pht_1_19 : _GEN_402; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_404 = 7'h14 == p1Addr ? pht_1_20 : _GEN_403; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_405 = 7'h15 == p1Addr ? pht_1_21 : _GEN_404; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_406 = 7'h16 == p1Addr ? pht_1_22 : _GEN_405; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_407 = 7'h17 == p1Addr ? pht_1_23 : _GEN_406; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_408 = 7'h18 == p1Addr ? pht_1_24 : _GEN_407; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_409 = 7'h19 == p1Addr ? pht_1_25 : _GEN_408; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_410 = 7'h1a == p1Addr ? pht_1_26 : _GEN_409; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_411 = 7'h1b == p1Addr ? pht_1_27 : _GEN_410; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_412 = 7'h1c == p1Addr ? pht_1_28 : _GEN_411; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_413 = 7'h1d == p1Addr ? pht_1_29 : _GEN_412; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_414 = 7'h1e == p1Addr ? pht_1_30 : _GEN_413; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_415 = 7'h1f == p1Addr ? pht_1_31 : _GEN_414; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_416 = 7'h20 == p1Addr ? pht_1_32 : _GEN_415; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_417 = 7'h21 == p1Addr ? pht_1_33 : _GEN_416; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_418 = 7'h22 == p1Addr ? pht_1_34 : _GEN_417; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_419 = 7'h23 == p1Addr ? pht_1_35 : _GEN_418; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_420 = 7'h24 == p1Addr ? pht_1_36 : _GEN_419; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_421 = 7'h25 == p1Addr ? pht_1_37 : _GEN_420; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_422 = 7'h26 == p1Addr ? pht_1_38 : _GEN_421; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_423 = 7'h27 == p1Addr ? pht_1_39 : _GEN_422; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_424 = 7'h28 == p1Addr ? pht_1_40 : _GEN_423; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_425 = 7'h29 == p1Addr ? pht_1_41 : _GEN_424; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_426 = 7'h2a == p1Addr ? pht_1_42 : _GEN_425; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_427 = 7'h2b == p1Addr ? pht_1_43 : _GEN_426; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_428 = 7'h2c == p1Addr ? pht_1_44 : _GEN_427; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_429 = 7'h2d == p1Addr ? pht_1_45 : _GEN_428; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_430 = 7'h2e == p1Addr ? pht_1_46 : _GEN_429; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_431 = 7'h2f == p1Addr ? pht_1_47 : _GEN_430; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_432 = 7'h30 == p1Addr ? pht_1_48 : _GEN_431; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_433 = 7'h31 == p1Addr ? pht_1_49 : _GEN_432; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_434 = 7'h32 == p1Addr ? pht_1_50 : _GEN_433; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_435 = 7'h33 == p1Addr ? pht_1_51 : _GEN_434; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_436 = 7'h34 == p1Addr ? pht_1_52 : _GEN_435; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_437 = 7'h35 == p1Addr ? pht_1_53 : _GEN_436; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_438 = 7'h36 == p1Addr ? pht_1_54 : _GEN_437; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_439 = 7'h37 == p1Addr ? pht_1_55 : _GEN_438; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_440 = 7'h38 == p1Addr ? pht_1_56 : _GEN_439; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_441 = 7'h39 == p1Addr ? pht_1_57 : _GEN_440; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_442 = 7'h3a == p1Addr ? pht_1_58 : _GEN_441; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_443 = 7'h3b == p1Addr ? pht_1_59 : _GEN_442; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_444 = 7'h3c == p1Addr ? pht_1_60 : _GEN_443; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_445 = 7'h3d == p1Addr ? pht_1_61 : _GEN_444; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_446 = 7'h3e == p1Addr ? pht_1_62 : _GEN_445; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_447 = 7'h3f == p1Addr ? pht_1_63 : _GEN_446; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_448 = 7'h40 == p1Addr ? pht_1_64 : _GEN_447; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_449 = 7'h41 == p1Addr ? pht_1_65 : _GEN_448; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_450 = 7'h42 == p1Addr ? pht_1_66 : _GEN_449; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_451 = 7'h43 == p1Addr ? pht_1_67 : _GEN_450; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_452 = 7'h44 == p1Addr ? pht_1_68 : _GEN_451; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_453 = 7'h45 == p1Addr ? pht_1_69 : _GEN_452; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_454 = 7'h46 == p1Addr ? pht_1_70 : _GEN_453; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_455 = 7'h47 == p1Addr ? pht_1_71 : _GEN_454; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_456 = 7'h48 == p1Addr ? pht_1_72 : _GEN_455; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_457 = 7'h49 == p1Addr ? pht_1_73 : _GEN_456; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_458 = 7'h4a == p1Addr ? pht_1_74 : _GEN_457; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_459 = 7'h4b == p1Addr ? pht_1_75 : _GEN_458; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_460 = 7'h4c == p1Addr ? pht_1_76 : _GEN_459; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_461 = 7'h4d == p1Addr ? pht_1_77 : _GEN_460; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_462 = 7'h4e == p1Addr ? pht_1_78 : _GEN_461; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_463 = 7'h4f == p1Addr ? pht_1_79 : _GEN_462; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_464 = 7'h50 == p1Addr ? pht_1_80 : _GEN_463; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_465 = 7'h51 == p1Addr ? pht_1_81 : _GEN_464; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_466 = 7'h52 == p1Addr ? pht_1_82 : _GEN_465; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_467 = 7'h53 == p1Addr ? pht_1_83 : _GEN_466; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_468 = 7'h54 == p1Addr ? pht_1_84 : _GEN_467; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_469 = 7'h55 == p1Addr ? pht_1_85 : _GEN_468; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_470 = 7'h56 == p1Addr ? pht_1_86 : _GEN_469; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_471 = 7'h57 == p1Addr ? pht_1_87 : _GEN_470; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_472 = 7'h58 == p1Addr ? pht_1_88 : _GEN_471; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_473 = 7'h59 == p1Addr ? pht_1_89 : _GEN_472; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_474 = 7'h5a == p1Addr ? pht_1_90 : _GEN_473; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_475 = 7'h5b == p1Addr ? pht_1_91 : _GEN_474; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_476 = 7'h5c == p1Addr ? pht_1_92 : _GEN_475; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_477 = 7'h5d == p1Addr ? pht_1_93 : _GEN_476; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_478 = 7'h5e == p1Addr ? pht_1_94 : _GEN_477; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_479 = 7'h5f == p1Addr ? pht_1_95 : _GEN_478; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_480 = 7'h60 == p1Addr ? pht_1_96 : _GEN_479; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_481 = 7'h61 == p1Addr ? pht_1_97 : _GEN_480; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_482 = 7'h62 == p1Addr ? pht_1_98 : _GEN_481; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_483 = 7'h63 == p1Addr ? pht_1_99 : _GEN_482; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_484 = 7'h64 == p1Addr ? pht_1_100 : _GEN_483; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_485 = 7'h65 == p1Addr ? pht_1_101 : _GEN_484; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_486 = 7'h66 == p1Addr ? pht_1_102 : _GEN_485; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_487 = 7'h67 == p1Addr ? pht_1_103 : _GEN_486; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_488 = 7'h68 == p1Addr ? pht_1_104 : _GEN_487; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_489 = 7'h69 == p1Addr ? pht_1_105 : _GEN_488; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_490 = 7'h6a == p1Addr ? pht_1_106 : _GEN_489; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_491 = 7'h6b == p1Addr ? pht_1_107 : _GEN_490; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_492 = 7'h6c == p1Addr ? pht_1_108 : _GEN_491; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_493 = 7'h6d == p1Addr ? pht_1_109 : _GEN_492; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_494 = 7'h6e == p1Addr ? pht_1_110 : _GEN_493; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_495 = 7'h6f == p1Addr ? pht_1_111 : _GEN_494; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_496 = 7'h70 == p1Addr ? pht_1_112 : _GEN_495; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_497 = 7'h71 == p1Addr ? pht_1_113 : _GEN_496; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_498 = 7'h72 == p1Addr ? pht_1_114 : _GEN_497; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_499 = 7'h73 == p1Addr ? pht_1_115 : _GEN_498; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_500 = 7'h74 == p1Addr ? pht_1_116 : _GEN_499; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_501 = 7'h75 == p1Addr ? pht_1_117 : _GEN_500; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_502 = 7'h76 == p1Addr ? pht_1_118 : _GEN_501; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_503 = 7'h77 == p1Addr ? pht_1_119 : _GEN_502; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_504 = 7'h78 == p1Addr ? pht_1_120 : _GEN_503; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_505 = 7'h79 == p1Addr ? pht_1_121 : _GEN_504; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_506 = 7'h7a == p1Addr ? pht_1_122 : _GEN_505; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_507 = 7'h7b == p1Addr ? pht_1_123 : _GEN_506; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_508 = 7'h7c == p1Addr ? pht_1_124 : _GEN_507; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_509 = 7'h7d == p1Addr ? pht_1_125 : _GEN_508; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_510 = 7'h7e == p1Addr ? pht_1_126 : _GEN_509; // @[bht.scala 123:{23,23}]
  wire [1:0] _GEN_511 = 7'h7f == p1Addr ? pht_1_127 : _GEN_510; // @[bht.scala 123:{23,23}]
  wire [1:0] phtData = _GEN_255[1] ? _GEN_383 : _GEN_511; // @[bht.scala 123:23]
  wire [6:0] reqIndex = io_pc[10:4]; // @[bht.scala 127:25]
  wire  _GEN_513 = 7'h1 == reqIndex ? btbV_1 : btbV_0; // @[bht.scala 128:{53,53}]
  wire  _GEN_514 = 7'h2 == reqIndex ? btbV_2 : _GEN_513; // @[bht.scala 128:{53,53}]
  wire  _GEN_515 = 7'h3 == reqIndex ? btbV_3 : _GEN_514; // @[bht.scala 128:{53,53}]
  wire  _GEN_516 = 7'h4 == reqIndex ? btbV_4 : _GEN_515; // @[bht.scala 128:{53,53}]
  wire  _GEN_517 = 7'h5 == reqIndex ? btbV_5 : _GEN_516; // @[bht.scala 128:{53,53}]
  wire  _GEN_518 = 7'h6 == reqIndex ? btbV_6 : _GEN_517; // @[bht.scala 128:{53,53}]
  wire  _GEN_519 = 7'h7 == reqIndex ? btbV_7 : _GEN_518; // @[bht.scala 128:{53,53}]
  wire  _GEN_520 = 7'h8 == reqIndex ? btbV_8 : _GEN_519; // @[bht.scala 128:{53,53}]
  wire  _GEN_521 = 7'h9 == reqIndex ? btbV_9 : _GEN_520; // @[bht.scala 128:{53,53}]
  wire  _GEN_522 = 7'ha == reqIndex ? btbV_10 : _GEN_521; // @[bht.scala 128:{53,53}]
  wire  _GEN_523 = 7'hb == reqIndex ? btbV_11 : _GEN_522; // @[bht.scala 128:{53,53}]
  wire  _GEN_524 = 7'hc == reqIndex ? btbV_12 : _GEN_523; // @[bht.scala 128:{53,53}]
  wire  _GEN_525 = 7'hd == reqIndex ? btbV_13 : _GEN_524; // @[bht.scala 128:{53,53}]
  wire  _GEN_526 = 7'he == reqIndex ? btbV_14 : _GEN_525; // @[bht.scala 128:{53,53}]
  wire  _GEN_527 = 7'hf == reqIndex ? btbV_15 : _GEN_526; // @[bht.scala 128:{53,53}]
  wire  _GEN_528 = 7'h10 == reqIndex ? btbV_16 : _GEN_527; // @[bht.scala 128:{53,53}]
  wire  _GEN_529 = 7'h11 == reqIndex ? btbV_17 : _GEN_528; // @[bht.scala 128:{53,53}]
  wire  _GEN_530 = 7'h12 == reqIndex ? btbV_18 : _GEN_529; // @[bht.scala 128:{53,53}]
  wire  _GEN_531 = 7'h13 == reqIndex ? btbV_19 : _GEN_530; // @[bht.scala 128:{53,53}]
  wire  _GEN_532 = 7'h14 == reqIndex ? btbV_20 : _GEN_531; // @[bht.scala 128:{53,53}]
  wire  _GEN_533 = 7'h15 == reqIndex ? btbV_21 : _GEN_532; // @[bht.scala 128:{53,53}]
  wire  _GEN_534 = 7'h16 == reqIndex ? btbV_22 : _GEN_533; // @[bht.scala 128:{53,53}]
  wire  _GEN_535 = 7'h17 == reqIndex ? btbV_23 : _GEN_534; // @[bht.scala 128:{53,53}]
  wire  _GEN_536 = 7'h18 == reqIndex ? btbV_24 : _GEN_535; // @[bht.scala 128:{53,53}]
  wire  _GEN_537 = 7'h19 == reqIndex ? btbV_25 : _GEN_536; // @[bht.scala 128:{53,53}]
  wire  _GEN_538 = 7'h1a == reqIndex ? btbV_26 : _GEN_537; // @[bht.scala 128:{53,53}]
  wire  _GEN_539 = 7'h1b == reqIndex ? btbV_27 : _GEN_538; // @[bht.scala 128:{53,53}]
  wire  _GEN_540 = 7'h1c == reqIndex ? btbV_28 : _GEN_539; // @[bht.scala 128:{53,53}]
  wire  _GEN_541 = 7'h1d == reqIndex ? btbV_29 : _GEN_540; // @[bht.scala 128:{53,53}]
  wire  _GEN_542 = 7'h1e == reqIndex ? btbV_30 : _GEN_541; // @[bht.scala 128:{53,53}]
  wire  _GEN_543 = 7'h1f == reqIndex ? btbV_31 : _GEN_542; // @[bht.scala 128:{53,53}]
  wire  _GEN_544 = 7'h20 == reqIndex ? btbV_32 : _GEN_543; // @[bht.scala 128:{53,53}]
  wire  _GEN_545 = 7'h21 == reqIndex ? btbV_33 : _GEN_544; // @[bht.scala 128:{53,53}]
  wire  _GEN_546 = 7'h22 == reqIndex ? btbV_34 : _GEN_545; // @[bht.scala 128:{53,53}]
  wire  _GEN_547 = 7'h23 == reqIndex ? btbV_35 : _GEN_546; // @[bht.scala 128:{53,53}]
  wire  _GEN_548 = 7'h24 == reqIndex ? btbV_36 : _GEN_547; // @[bht.scala 128:{53,53}]
  wire  _GEN_549 = 7'h25 == reqIndex ? btbV_37 : _GEN_548; // @[bht.scala 128:{53,53}]
  wire  _GEN_550 = 7'h26 == reqIndex ? btbV_38 : _GEN_549; // @[bht.scala 128:{53,53}]
  wire  _GEN_551 = 7'h27 == reqIndex ? btbV_39 : _GEN_550; // @[bht.scala 128:{53,53}]
  wire  _GEN_552 = 7'h28 == reqIndex ? btbV_40 : _GEN_551; // @[bht.scala 128:{53,53}]
  wire  _GEN_553 = 7'h29 == reqIndex ? btbV_41 : _GEN_552; // @[bht.scala 128:{53,53}]
  wire  _GEN_554 = 7'h2a == reqIndex ? btbV_42 : _GEN_553; // @[bht.scala 128:{53,53}]
  wire  _GEN_555 = 7'h2b == reqIndex ? btbV_43 : _GEN_554; // @[bht.scala 128:{53,53}]
  wire  _GEN_556 = 7'h2c == reqIndex ? btbV_44 : _GEN_555; // @[bht.scala 128:{53,53}]
  wire  _GEN_557 = 7'h2d == reqIndex ? btbV_45 : _GEN_556; // @[bht.scala 128:{53,53}]
  wire  _GEN_558 = 7'h2e == reqIndex ? btbV_46 : _GEN_557; // @[bht.scala 128:{53,53}]
  wire  _GEN_559 = 7'h2f == reqIndex ? btbV_47 : _GEN_558; // @[bht.scala 128:{53,53}]
  wire  _GEN_560 = 7'h30 == reqIndex ? btbV_48 : _GEN_559; // @[bht.scala 128:{53,53}]
  wire  _GEN_561 = 7'h31 == reqIndex ? btbV_49 : _GEN_560; // @[bht.scala 128:{53,53}]
  wire  _GEN_562 = 7'h32 == reqIndex ? btbV_50 : _GEN_561; // @[bht.scala 128:{53,53}]
  wire  _GEN_563 = 7'h33 == reqIndex ? btbV_51 : _GEN_562; // @[bht.scala 128:{53,53}]
  wire  _GEN_564 = 7'h34 == reqIndex ? btbV_52 : _GEN_563; // @[bht.scala 128:{53,53}]
  wire  _GEN_565 = 7'h35 == reqIndex ? btbV_53 : _GEN_564; // @[bht.scala 128:{53,53}]
  wire  _GEN_566 = 7'h36 == reqIndex ? btbV_54 : _GEN_565; // @[bht.scala 128:{53,53}]
  wire  _GEN_567 = 7'h37 == reqIndex ? btbV_55 : _GEN_566; // @[bht.scala 128:{53,53}]
  wire  _GEN_568 = 7'h38 == reqIndex ? btbV_56 : _GEN_567; // @[bht.scala 128:{53,53}]
  wire  _GEN_569 = 7'h39 == reqIndex ? btbV_57 : _GEN_568; // @[bht.scala 128:{53,53}]
  wire  _GEN_570 = 7'h3a == reqIndex ? btbV_58 : _GEN_569; // @[bht.scala 128:{53,53}]
  wire  _GEN_571 = 7'h3b == reqIndex ? btbV_59 : _GEN_570; // @[bht.scala 128:{53,53}]
  wire  _GEN_572 = 7'h3c == reqIndex ? btbV_60 : _GEN_571; // @[bht.scala 128:{53,53}]
  wire  _GEN_573 = 7'h3d == reqIndex ? btbV_61 : _GEN_572; // @[bht.scala 128:{53,53}]
  wire  _GEN_574 = 7'h3e == reqIndex ? btbV_62 : _GEN_573; // @[bht.scala 128:{53,53}]
  wire  _GEN_575 = 7'h3f == reqIndex ? btbV_63 : _GEN_574; // @[bht.scala 128:{53,53}]
  wire  _GEN_576 = 7'h40 == reqIndex ? btbV_64 : _GEN_575; // @[bht.scala 128:{53,53}]
  wire  _GEN_577 = 7'h41 == reqIndex ? btbV_65 : _GEN_576; // @[bht.scala 128:{53,53}]
  wire  _GEN_578 = 7'h42 == reqIndex ? btbV_66 : _GEN_577; // @[bht.scala 128:{53,53}]
  wire  _GEN_579 = 7'h43 == reqIndex ? btbV_67 : _GEN_578; // @[bht.scala 128:{53,53}]
  wire  _GEN_580 = 7'h44 == reqIndex ? btbV_68 : _GEN_579; // @[bht.scala 128:{53,53}]
  wire  _GEN_581 = 7'h45 == reqIndex ? btbV_69 : _GEN_580; // @[bht.scala 128:{53,53}]
  wire  _GEN_582 = 7'h46 == reqIndex ? btbV_70 : _GEN_581; // @[bht.scala 128:{53,53}]
  wire  _GEN_583 = 7'h47 == reqIndex ? btbV_71 : _GEN_582; // @[bht.scala 128:{53,53}]
  wire  _GEN_584 = 7'h48 == reqIndex ? btbV_72 : _GEN_583; // @[bht.scala 128:{53,53}]
  wire  _GEN_585 = 7'h49 == reqIndex ? btbV_73 : _GEN_584; // @[bht.scala 128:{53,53}]
  wire  _GEN_586 = 7'h4a == reqIndex ? btbV_74 : _GEN_585; // @[bht.scala 128:{53,53}]
  wire  _GEN_587 = 7'h4b == reqIndex ? btbV_75 : _GEN_586; // @[bht.scala 128:{53,53}]
  wire  _GEN_588 = 7'h4c == reqIndex ? btbV_76 : _GEN_587; // @[bht.scala 128:{53,53}]
  wire  _GEN_589 = 7'h4d == reqIndex ? btbV_77 : _GEN_588; // @[bht.scala 128:{53,53}]
  wire  _GEN_590 = 7'h4e == reqIndex ? btbV_78 : _GEN_589; // @[bht.scala 128:{53,53}]
  wire  _GEN_591 = 7'h4f == reqIndex ? btbV_79 : _GEN_590; // @[bht.scala 128:{53,53}]
  wire  _GEN_592 = 7'h50 == reqIndex ? btbV_80 : _GEN_591; // @[bht.scala 128:{53,53}]
  wire  _GEN_593 = 7'h51 == reqIndex ? btbV_81 : _GEN_592; // @[bht.scala 128:{53,53}]
  wire  _GEN_594 = 7'h52 == reqIndex ? btbV_82 : _GEN_593; // @[bht.scala 128:{53,53}]
  wire  _GEN_595 = 7'h53 == reqIndex ? btbV_83 : _GEN_594; // @[bht.scala 128:{53,53}]
  wire  _GEN_596 = 7'h54 == reqIndex ? btbV_84 : _GEN_595; // @[bht.scala 128:{53,53}]
  wire  _GEN_597 = 7'h55 == reqIndex ? btbV_85 : _GEN_596; // @[bht.scala 128:{53,53}]
  wire  _GEN_598 = 7'h56 == reqIndex ? btbV_86 : _GEN_597; // @[bht.scala 128:{53,53}]
  wire  _GEN_599 = 7'h57 == reqIndex ? btbV_87 : _GEN_598; // @[bht.scala 128:{53,53}]
  wire  _GEN_600 = 7'h58 == reqIndex ? btbV_88 : _GEN_599; // @[bht.scala 128:{53,53}]
  wire  _GEN_601 = 7'h59 == reqIndex ? btbV_89 : _GEN_600; // @[bht.scala 128:{53,53}]
  wire  _GEN_602 = 7'h5a == reqIndex ? btbV_90 : _GEN_601; // @[bht.scala 128:{53,53}]
  wire  _GEN_603 = 7'h5b == reqIndex ? btbV_91 : _GEN_602; // @[bht.scala 128:{53,53}]
  wire  _GEN_604 = 7'h5c == reqIndex ? btbV_92 : _GEN_603; // @[bht.scala 128:{53,53}]
  wire  _GEN_605 = 7'h5d == reqIndex ? btbV_93 : _GEN_604; // @[bht.scala 128:{53,53}]
  wire  _GEN_606 = 7'h5e == reqIndex ? btbV_94 : _GEN_605; // @[bht.scala 128:{53,53}]
  wire  _GEN_607 = 7'h5f == reqIndex ? btbV_95 : _GEN_606; // @[bht.scala 128:{53,53}]
  wire  _GEN_608 = 7'h60 == reqIndex ? btbV_96 : _GEN_607; // @[bht.scala 128:{53,53}]
  wire  _GEN_609 = 7'h61 == reqIndex ? btbV_97 : _GEN_608; // @[bht.scala 128:{53,53}]
  wire  _GEN_610 = 7'h62 == reqIndex ? btbV_98 : _GEN_609; // @[bht.scala 128:{53,53}]
  wire  _GEN_611 = 7'h63 == reqIndex ? btbV_99 : _GEN_610; // @[bht.scala 128:{53,53}]
  wire  _GEN_612 = 7'h64 == reqIndex ? btbV_100 : _GEN_611; // @[bht.scala 128:{53,53}]
  wire  _GEN_613 = 7'h65 == reqIndex ? btbV_101 : _GEN_612; // @[bht.scala 128:{53,53}]
  wire  _GEN_614 = 7'h66 == reqIndex ? btbV_102 : _GEN_613; // @[bht.scala 128:{53,53}]
  wire  _GEN_615 = 7'h67 == reqIndex ? btbV_103 : _GEN_614; // @[bht.scala 128:{53,53}]
  wire  _GEN_616 = 7'h68 == reqIndex ? btbV_104 : _GEN_615; // @[bht.scala 128:{53,53}]
  wire  _GEN_617 = 7'h69 == reqIndex ? btbV_105 : _GEN_616; // @[bht.scala 128:{53,53}]
  wire  _GEN_618 = 7'h6a == reqIndex ? btbV_106 : _GEN_617; // @[bht.scala 128:{53,53}]
  wire  _GEN_619 = 7'h6b == reqIndex ? btbV_107 : _GEN_618; // @[bht.scala 128:{53,53}]
  wire  _GEN_620 = 7'h6c == reqIndex ? btbV_108 : _GEN_619; // @[bht.scala 128:{53,53}]
  wire  _GEN_621 = 7'h6d == reqIndex ? btbV_109 : _GEN_620; // @[bht.scala 128:{53,53}]
  wire  _GEN_622 = 7'h6e == reqIndex ? btbV_110 : _GEN_621; // @[bht.scala 128:{53,53}]
  wire  _GEN_623 = 7'h6f == reqIndex ? btbV_111 : _GEN_622; // @[bht.scala 128:{53,53}]
  wire  _GEN_624 = 7'h70 == reqIndex ? btbV_112 : _GEN_623; // @[bht.scala 128:{53,53}]
  wire  _GEN_625 = 7'h71 == reqIndex ? btbV_113 : _GEN_624; // @[bht.scala 128:{53,53}]
  wire  _GEN_626 = 7'h72 == reqIndex ? btbV_114 : _GEN_625; // @[bht.scala 128:{53,53}]
  wire  _GEN_627 = 7'h73 == reqIndex ? btbV_115 : _GEN_626; // @[bht.scala 128:{53,53}]
  wire  _GEN_628 = 7'h74 == reqIndex ? btbV_116 : _GEN_627; // @[bht.scala 128:{53,53}]
  wire  _GEN_629 = 7'h75 == reqIndex ? btbV_117 : _GEN_628; // @[bht.scala 128:{53,53}]
  wire  _GEN_630 = 7'h76 == reqIndex ? btbV_118 : _GEN_629; // @[bht.scala 128:{53,53}]
  wire  _GEN_631 = 7'h77 == reqIndex ? btbV_119 : _GEN_630; // @[bht.scala 128:{53,53}]
  wire  _GEN_632 = 7'h78 == reqIndex ? btbV_120 : _GEN_631; // @[bht.scala 128:{53,53}]
  wire  _GEN_633 = 7'h79 == reqIndex ? btbV_121 : _GEN_632; // @[bht.scala 128:{53,53}]
  wire  _GEN_634 = 7'h7a == reqIndex ? btbV_122 : _GEN_633; // @[bht.scala 128:{53,53}]
  wire  _GEN_635 = 7'h7b == reqIndex ? btbV_123 : _GEN_634; // @[bht.scala 128:{53,53}]
  wire  _GEN_636 = 7'h7c == reqIndex ? btbV_124 : _GEN_635; // @[bht.scala 128:{53,53}]
  wire  _GEN_637 = 7'h7d == reqIndex ? btbV_125 : _GEN_636; // @[bht.scala 128:{53,53}]
  wire  _GEN_638 = 7'h7e == reqIndex ? btbV_126 : _GEN_637; // @[bht.scala 128:{53,53}]
  wire  _GEN_639 = 7'h7f == reqIndex ? btbV_127 : _GEN_638; // @[bht.scala 128:{53,53}]
  wire [6:0] _GEN_641 = 7'h1 == reqIndex ? btbTag_1 : btbTag_0; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_642 = 7'h2 == reqIndex ? btbTag_2 : _GEN_641; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_643 = 7'h3 == reqIndex ? btbTag_3 : _GEN_642; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_644 = 7'h4 == reqIndex ? btbTag_4 : _GEN_643; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_645 = 7'h5 == reqIndex ? btbTag_5 : _GEN_644; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_646 = 7'h6 == reqIndex ? btbTag_6 : _GEN_645; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_647 = 7'h7 == reqIndex ? btbTag_7 : _GEN_646; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_648 = 7'h8 == reqIndex ? btbTag_8 : _GEN_647; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_649 = 7'h9 == reqIndex ? btbTag_9 : _GEN_648; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_650 = 7'ha == reqIndex ? btbTag_10 : _GEN_649; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_651 = 7'hb == reqIndex ? btbTag_11 : _GEN_650; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_652 = 7'hc == reqIndex ? btbTag_12 : _GEN_651; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_653 = 7'hd == reqIndex ? btbTag_13 : _GEN_652; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_654 = 7'he == reqIndex ? btbTag_14 : _GEN_653; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_655 = 7'hf == reqIndex ? btbTag_15 : _GEN_654; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_656 = 7'h10 == reqIndex ? btbTag_16 : _GEN_655; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_657 = 7'h11 == reqIndex ? btbTag_17 : _GEN_656; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_658 = 7'h12 == reqIndex ? btbTag_18 : _GEN_657; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_659 = 7'h13 == reqIndex ? btbTag_19 : _GEN_658; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_660 = 7'h14 == reqIndex ? btbTag_20 : _GEN_659; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_661 = 7'h15 == reqIndex ? btbTag_21 : _GEN_660; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_662 = 7'h16 == reqIndex ? btbTag_22 : _GEN_661; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_663 = 7'h17 == reqIndex ? btbTag_23 : _GEN_662; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_664 = 7'h18 == reqIndex ? btbTag_24 : _GEN_663; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_665 = 7'h19 == reqIndex ? btbTag_25 : _GEN_664; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_666 = 7'h1a == reqIndex ? btbTag_26 : _GEN_665; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_667 = 7'h1b == reqIndex ? btbTag_27 : _GEN_666; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_668 = 7'h1c == reqIndex ? btbTag_28 : _GEN_667; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_669 = 7'h1d == reqIndex ? btbTag_29 : _GEN_668; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_670 = 7'h1e == reqIndex ? btbTag_30 : _GEN_669; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_671 = 7'h1f == reqIndex ? btbTag_31 : _GEN_670; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_672 = 7'h20 == reqIndex ? btbTag_32 : _GEN_671; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_673 = 7'h21 == reqIndex ? btbTag_33 : _GEN_672; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_674 = 7'h22 == reqIndex ? btbTag_34 : _GEN_673; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_675 = 7'h23 == reqIndex ? btbTag_35 : _GEN_674; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_676 = 7'h24 == reqIndex ? btbTag_36 : _GEN_675; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_677 = 7'h25 == reqIndex ? btbTag_37 : _GEN_676; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_678 = 7'h26 == reqIndex ? btbTag_38 : _GEN_677; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_679 = 7'h27 == reqIndex ? btbTag_39 : _GEN_678; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_680 = 7'h28 == reqIndex ? btbTag_40 : _GEN_679; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_681 = 7'h29 == reqIndex ? btbTag_41 : _GEN_680; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_682 = 7'h2a == reqIndex ? btbTag_42 : _GEN_681; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_683 = 7'h2b == reqIndex ? btbTag_43 : _GEN_682; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_684 = 7'h2c == reqIndex ? btbTag_44 : _GEN_683; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_685 = 7'h2d == reqIndex ? btbTag_45 : _GEN_684; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_686 = 7'h2e == reqIndex ? btbTag_46 : _GEN_685; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_687 = 7'h2f == reqIndex ? btbTag_47 : _GEN_686; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_688 = 7'h30 == reqIndex ? btbTag_48 : _GEN_687; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_689 = 7'h31 == reqIndex ? btbTag_49 : _GEN_688; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_690 = 7'h32 == reqIndex ? btbTag_50 : _GEN_689; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_691 = 7'h33 == reqIndex ? btbTag_51 : _GEN_690; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_692 = 7'h34 == reqIndex ? btbTag_52 : _GEN_691; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_693 = 7'h35 == reqIndex ? btbTag_53 : _GEN_692; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_694 = 7'h36 == reqIndex ? btbTag_54 : _GEN_693; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_695 = 7'h37 == reqIndex ? btbTag_55 : _GEN_694; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_696 = 7'h38 == reqIndex ? btbTag_56 : _GEN_695; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_697 = 7'h39 == reqIndex ? btbTag_57 : _GEN_696; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_698 = 7'h3a == reqIndex ? btbTag_58 : _GEN_697; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_699 = 7'h3b == reqIndex ? btbTag_59 : _GEN_698; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_700 = 7'h3c == reqIndex ? btbTag_60 : _GEN_699; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_701 = 7'h3d == reqIndex ? btbTag_61 : _GEN_700; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_702 = 7'h3e == reqIndex ? btbTag_62 : _GEN_701; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_703 = 7'h3f == reqIndex ? btbTag_63 : _GEN_702; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_704 = 7'h40 == reqIndex ? btbTag_64 : _GEN_703; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_705 = 7'h41 == reqIndex ? btbTag_65 : _GEN_704; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_706 = 7'h42 == reqIndex ? btbTag_66 : _GEN_705; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_707 = 7'h43 == reqIndex ? btbTag_67 : _GEN_706; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_708 = 7'h44 == reqIndex ? btbTag_68 : _GEN_707; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_709 = 7'h45 == reqIndex ? btbTag_69 : _GEN_708; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_710 = 7'h46 == reqIndex ? btbTag_70 : _GEN_709; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_711 = 7'h47 == reqIndex ? btbTag_71 : _GEN_710; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_712 = 7'h48 == reqIndex ? btbTag_72 : _GEN_711; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_713 = 7'h49 == reqIndex ? btbTag_73 : _GEN_712; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_714 = 7'h4a == reqIndex ? btbTag_74 : _GEN_713; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_715 = 7'h4b == reqIndex ? btbTag_75 : _GEN_714; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_716 = 7'h4c == reqIndex ? btbTag_76 : _GEN_715; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_717 = 7'h4d == reqIndex ? btbTag_77 : _GEN_716; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_718 = 7'h4e == reqIndex ? btbTag_78 : _GEN_717; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_719 = 7'h4f == reqIndex ? btbTag_79 : _GEN_718; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_720 = 7'h50 == reqIndex ? btbTag_80 : _GEN_719; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_721 = 7'h51 == reqIndex ? btbTag_81 : _GEN_720; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_722 = 7'h52 == reqIndex ? btbTag_82 : _GEN_721; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_723 = 7'h53 == reqIndex ? btbTag_83 : _GEN_722; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_724 = 7'h54 == reqIndex ? btbTag_84 : _GEN_723; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_725 = 7'h55 == reqIndex ? btbTag_85 : _GEN_724; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_726 = 7'h56 == reqIndex ? btbTag_86 : _GEN_725; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_727 = 7'h57 == reqIndex ? btbTag_87 : _GEN_726; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_728 = 7'h58 == reqIndex ? btbTag_88 : _GEN_727; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_729 = 7'h59 == reqIndex ? btbTag_89 : _GEN_728; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_730 = 7'h5a == reqIndex ? btbTag_90 : _GEN_729; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_731 = 7'h5b == reqIndex ? btbTag_91 : _GEN_730; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_732 = 7'h5c == reqIndex ? btbTag_92 : _GEN_731; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_733 = 7'h5d == reqIndex ? btbTag_93 : _GEN_732; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_734 = 7'h5e == reqIndex ? btbTag_94 : _GEN_733; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_735 = 7'h5f == reqIndex ? btbTag_95 : _GEN_734; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_736 = 7'h60 == reqIndex ? btbTag_96 : _GEN_735; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_737 = 7'h61 == reqIndex ? btbTag_97 : _GEN_736; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_738 = 7'h62 == reqIndex ? btbTag_98 : _GEN_737; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_739 = 7'h63 == reqIndex ? btbTag_99 : _GEN_738; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_740 = 7'h64 == reqIndex ? btbTag_100 : _GEN_739; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_741 = 7'h65 == reqIndex ? btbTag_101 : _GEN_740; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_742 = 7'h66 == reqIndex ? btbTag_102 : _GEN_741; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_743 = 7'h67 == reqIndex ? btbTag_103 : _GEN_742; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_744 = 7'h68 == reqIndex ? btbTag_104 : _GEN_743; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_745 = 7'h69 == reqIndex ? btbTag_105 : _GEN_744; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_746 = 7'h6a == reqIndex ? btbTag_106 : _GEN_745; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_747 = 7'h6b == reqIndex ? btbTag_107 : _GEN_746; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_748 = 7'h6c == reqIndex ? btbTag_108 : _GEN_747; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_749 = 7'h6d == reqIndex ? btbTag_109 : _GEN_748; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_750 = 7'h6e == reqIndex ? btbTag_110 : _GEN_749; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_751 = 7'h6f == reqIndex ? btbTag_111 : _GEN_750; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_752 = 7'h70 == reqIndex ? btbTag_112 : _GEN_751; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_753 = 7'h71 == reqIndex ? btbTag_113 : _GEN_752; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_754 = 7'h72 == reqIndex ? btbTag_114 : _GEN_753; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_755 = 7'h73 == reqIndex ? btbTag_115 : _GEN_754; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_756 = 7'h74 == reqIndex ? btbTag_116 : _GEN_755; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_757 = 7'h75 == reqIndex ? btbTag_117 : _GEN_756; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_758 = 7'h76 == reqIndex ? btbTag_118 : _GEN_757; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_759 = 7'h77 == reqIndex ? btbTag_119 : _GEN_758; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_760 = 7'h78 == reqIndex ? btbTag_120 : _GEN_759; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_761 = 7'h79 == reqIndex ? btbTag_121 : _GEN_760; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_762 = 7'h7a == reqIndex ? btbTag_122 : _GEN_761; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_763 = 7'h7b == reqIndex ? btbTag_123 : _GEN_762; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_764 = 7'h7c == reqIndex ? btbTag_124 : _GEN_763; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_765 = 7'h7d == reqIndex ? btbTag_125 : _GEN_764; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_766 = 7'h7e == reqIndex ? btbTag_126 : _GEN_765; // @[bht.scala 128:{92,92}]
  wire [6:0] _GEN_767 = 7'h7f == reqIndex ? btbTag_127 : _GEN_766; // @[bht.scala 128:{92,92}]
  wire  btbHit = (io_bxx | io_jalr) & io_takenPre & _GEN_639 & _GEN_767 == _p1Addr_T_6; // @[bht.scala 128:71]
  wire  _io_takenPre_T_3 = io_bxx & phtData[1]; // @[bht.scala 134:26]
  wire  _io_takenPre_T_4 = io_jal | io_jalr | _io_takenPre_T_3; // @[bht.scala 133:24]
  wire [63:0] _io_takenPrePC_T_2 = op1 + io_imm; // @[bht.scala 138:47]
  wire [31:0] _GEN_769 = 7'h1 == reqIndex ? btbMeta_1 : btbMeta_0; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_770 = 7'h2 == reqIndex ? btbMeta_2 : _GEN_769; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_771 = 7'h3 == reqIndex ? btbMeta_3 : _GEN_770; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_772 = 7'h4 == reqIndex ? btbMeta_4 : _GEN_771; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_773 = 7'h5 == reqIndex ? btbMeta_5 : _GEN_772; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_774 = 7'h6 == reqIndex ? btbMeta_6 : _GEN_773; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_775 = 7'h7 == reqIndex ? btbMeta_7 : _GEN_774; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_776 = 7'h8 == reqIndex ? btbMeta_8 : _GEN_775; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_777 = 7'h9 == reqIndex ? btbMeta_9 : _GEN_776; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_778 = 7'ha == reqIndex ? btbMeta_10 : _GEN_777; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_779 = 7'hb == reqIndex ? btbMeta_11 : _GEN_778; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_780 = 7'hc == reqIndex ? btbMeta_12 : _GEN_779; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_781 = 7'hd == reqIndex ? btbMeta_13 : _GEN_780; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_782 = 7'he == reqIndex ? btbMeta_14 : _GEN_781; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_783 = 7'hf == reqIndex ? btbMeta_15 : _GEN_782; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_784 = 7'h10 == reqIndex ? btbMeta_16 : _GEN_783; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_785 = 7'h11 == reqIndex ? btbMeta_17 : _GEN_784; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_786 = 7'h12 == reqIndex ? btbMeta_18 : _GEN_785; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_787 = 7'h13 == reqIndex ? btbMeta_19 : _GEN_786; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_788 = 7'h14 == reqIndex ? btbMeta_20 : _GEN_787; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_789 = 7'h15 == reqIndex ? btbMeta_21 : _GEN_788; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_790 = 7'h16 == reqIndex ? btbMeta_22 : _GEN_789; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_791 = 7'h17 == reqIndex ? btbMeta_23 : _GEN_790; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_792 = 7'h18 == reqIndex ? btbMeta_24 : _GEN_791; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_793 = 7'h19 == reqIndex ? btbMeta_25 : _GEN_792; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_794 = 7'h1a == reqIndex ? btbMeta_26 : _GEN_793; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_795 = 7'h1b == reqIndex ? btbMeta_27 : _GEN_794; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_796 = 7'h1c == reqIndex ? btbMeta_28 : _GEN_795; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_797 = 7'h1d == reqIndex ? btbMeta_29 : _GEN_796; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_798 = 7'h1e == reqIndex ? btbMeta_30 : _GEN_797; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_799 = 7'h1f == reqIndex ? btbMeta_31 : _GEN_798; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_800 = 7'h20 == reqIndex ? btbMeta_32 : _GEN_799; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_801 = 7'h21 == reqIndex ? btbMeta_33 : _GEN_800; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_802 = 7'h22 == reqIndex ? btbMeta_34 : _GEN_801; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_803 = 7'h23 == reqIndex ? btbMeta_35 : _GEN_802; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_804 = 7'h24 == reqIndex ? btbMeta_36 : _GEN_803; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_805 = 7'h25 == reqIndex ? btbMeta_37 : _GEN_804; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_806 = 7'h26 == reqIndex ? btbMeta_38 : _GEN_805; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_807 = 7'h27 == reqIndex ? btbMeta_39 : _GEN_806; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_808 = 7'h28 == reqIndex ? btbMeta_40 : _GEN_807; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_809 = 7'h29 == reqIndex ? btbMeta_41 : _GEN_808; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_810 = 7'h2a == reqIndex ? btbMeta_42 : _GEN_809; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_811 = 7'h2b == reqIndex ? btbMeta_43 : _GEN_810; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_812 = 7'h2c == reqIndex ? btbMeta_44 : _GEN_811; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_813 = 7'h2d == reqIndex ? btbMeta_45 : _GEN_812; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_814 = 7'h2e == reqIndex ? btbMeta_46 : _GEN_813; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_815 = 7'h2f == reqIndex ? btbMeta_47 : _GEN_814; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_816 = 7'h30 == reqIndex ? btbMeta_48 : _GEN_815; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_817 = 7'h31 == reqIndex ? btbMeta_49 : _GEN_816; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_818 = 7'h32 == reqIndex ? btbMeta_50 : _GEN_817; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_819 = 7'h33 == reqIndex ? btbMeta_51 : _GEN_818; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_820 = 7'h34 == reqIndex ? btbMeta_52 : _GEN_819; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_821 = 7'h35 == reqIndex ? btbMeta_53 : _GEN_820; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_822 = 7'h36 == reqIndex ? btbMeta_54 : _GEN_821; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_823 = 7'h37 == reqIndex ? btbMeta_55 : _GEN_822; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_824 = 7'h38 == reqIndex ? btbMeta_56 : _GEN_823; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_825 = 7'h39 == reqIndex ? btbMeta_57 : _GEN_824; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_826 = 7'h3a == reqIndex ? btbMeta_58 : _GEN_825; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_827 = 7'h3b == reqIndex ? btbMeta_59 : _GEN_826; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_828 = 7'h3c == reqIndex ? btbMeta_60 : _GEN_827; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_829 = 7'h3d == reqIndex ? btbMeta_61 : _GEN_828; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_830 = 7'h3e == reqIndex ? btbMeta_62 : _GEN_829; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_831 = 7'h3f == reqIndex ? btbMeta_63 : _GEN_830; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_832 = 7'h40 == reqIndex ? btbMeta_64 : _GEN_831; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_833 = 7'h41 == reqIndex ? btbMeta_65 : _GEN_832; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_834 = 7'h42 == reqIndex ? btbMeta_66 : _GEN_833; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_835 = 7'h43 == reqIndex ? btbMeta_67 : _GEN_834; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_836 = 7'h44 == reqIndex ? btbMeta_68 : _GEN_835; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_837 = 7'h45 == reqIndex ? btbMeta_69 : _GEN_836; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_838 = 7'h46 == reqIndex ? btbMeta_70 : _GEN_837; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_839 = 7'h47 == reqIndex ? btbMeta_71 : _GEN_838; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_840 = 7'h48 == reqIndex ? btbMeta_72 : _GEN_839; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_841 = 7'h49 == reqIndex ? btbMeta_73 : _GEN_840; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_842 = 7'h4a == reqIndex ? btbMeta_74 : _GEN_841; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_843 = 7'h4b == reqIndex ? btbMeta_75 : _GEN_842; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_844 = 7'h4c == reqIndex ? btbMeta_76 : _GEN_843; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_845 = 7'h4d == reqIndex ? btbMeta_77 : _GEN_844; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_846 = 7'h4e == reqIndex ? btbMeta_78 : _GEN_845; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_847 = 7'h4f == reqIndex ? btbMeta_79 : _GEN_846; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_848 = 7'h50 == reqIndex ? btbMeta_80 : _GEN_847; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_849 = 7'h51 == reqIndex ? btbMeta_81 : _GEN_848; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_850 = 7'h52 == reqIndex ? btbMeta_82 : _GEN_849; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_851 = 7'h53 == reqIndex ? btbMeta_83 : _GEN_850; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_852 = 7'h54 == reqIndex ? btbMeta_84 : _GEN_851; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_853 = 7'h55 == reqIndex ? btbMeta_85 : _GEN_852; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_854 = 7'h56 == reqIndex ? btbMeta_86 : _GEN_853; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_855 = 7'h57 == reqIndex ? btbMeta_87 : _GEN_854; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_856 = 7'h58 == reqIndex ? btbMeta_88 : _GEN_855; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_857 = 7'h59 == reqIndex ? btbMeta_89 : _GEN_856; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_858 = 7'h5a == reqIndex ? btbMeta_90 : _GEN_857; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_859 = 7'h5b == reqIndex ? btbMeta_91 : _GEN_858; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_860 = 7'h5c == reqIndex ? btbMeta_92 : _GEN_859; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_861 = 7'h5d == reqIndex ? btbMeta_93 : _GEN_860; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_862 = 7'h5e == reqIndex ? btbMeta_94 : _GEN_861; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_863 = 7'h5f == reqIndex ? btbMeta_95 : _GEN_862; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_864 = 7'h60 == reqIndex ? btbMeta_96 : _GEN_863; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_865 = 7'h61 == reqIndex ? btbMeta_97 : _GEN_864; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_866 = 7'h62 == reqIndex ? btbMeta_98 : _GEN_865; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_867 = 7'h63 == reqIndex ? btbMeta_99 : _GEN_866; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_868 = 7'h64 == reqIndex ? btbMeta_100 : _GEN_867; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_869 = 7'h65 == reqIndex ? btbMeta_101 : _GEN_868; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_870 = 7'h66 == reqIndex ? btbMeta_102 : _GEN_869; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_871 = 7'h67 == reqIndex ? btbMeta_103 : _GEN_870; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_872 = 7'h68 == reqIndex ? btbMeta_104 : _GEN_871; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_873 = 7'h69 == reqIndex ? btbMeta_105 : _GEN_872; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_874 = 7'h6a == reqIndex ? btbMeta_106 : _GEN_873; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_875 = 7'h6b == reqIndex ? btbMeta_107 : _GEN_874; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_876 = 7'h6c == reqIndex ? btbMeta_108 : _GEN_875; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_877 = 7'h6d == reqIndex ? btbMeta_109 : _GEN_876; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_878 = 7'h6e == reqIndex ? btbMeta_110 : _GEN_877; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_879 = 7'h6f == reqIndex ? btbMeta_111 : _GEN_878; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_880 = 7'h70 == reqIndex ? btbMeta_112 : _GEN_879; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_881 = 7'h71 == reqIndex ? btbMeta_113 : _GEN_880; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_882 = 7'h72 == reqIndex ? btbMeta_114 : _GEN_881; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_883 = 7'h73 == reqIndex ? btbMeta_115 : _GEN_882; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_884 = 7'h74 == reqIndex ? btbMeta_116 : _GEN_883; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_885 = 7'h75 == reqIndex ? btbMeta_117 : _GEN_884; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_886 = 7'h76 == reqIndex ? btbMeta_118 : _GEN_885; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_887 = 7'h77 == reqIndex ? btbMeta_119 : _GEN_886; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_888 = 7'h78 == reqIndex ? btbMeta_120 : _GEN_887; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_889 = 7'h79 == reqIndex ? btbMeta_121 : _GEN_888; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_890 = 7'h7a == reqIndex ? btbMeta_122 : _GEN_889; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_891 = 7'h7b == reqIndex ? btbMeta_123 : _GEN_890; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_892 = 7'h7c == reqIndex ? btbMeta_124 : _GEN_891; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_893 = 7'h7d == reqIndex ? btbMeta_125 : _GEN_892; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_894 = 7'h7e == reqIndex ? btbMeta_126 : _GEN_893; // @[bht.scala 138:{26,26}]
  wire [31:0] _GEN_895 = 7'h7f == reqIndex ? btbMeta_127 : _GEN_894; // @[bht.scala 138:{26,26}]
  wire [63:0] _io_takenPrePC_T_3 = btbHit ? {{32'd0}, _GEN_895} : _io_takenPrePC_T_2; // @[bht.scala 138:26]
  wire [63:0] _io_takenPrePC_T_4 = io_valid & io_takenPre ? _io_takenPrePC_T_3 : 64'h0; // @[bht.scala 137:25]
  reg  io_ready_REG; // @[bht.scala 142:48]
  wire  bhtWAddr_hash0 = io_takenPC[2] ^ io_takenPC[14]; // @[bht.scala 90:27]
  wire  _bhtWAddr_hash1_T_2 = io_takenPC[9] ^ io_takenPC[10]; // @[bht.scala 91:28]
  wire  bhtWAddr_hash1 = io_takenPC[9] ^ io_takenPC[10] ^ (io_takenPC[3] ^ io_takenPC[15]); // @[bht.scala 91:39]
  wire  bhtWAddr_hash2 = io_takenPC[4] ^ (io_takenPC[10] ^ io_takenPC[11]); // @[bht.scala 92:27]
  wire  bhtWAddr_hash3 = io_takenPC[5] ^ (io_takenPC[11] ^ io_takenPC[12]); // @[bht.scala 93:27]
  wire  bhtWAddr_hash4 = io_takenPC[6] ^ (io_takenPC[12] ^ io_takenPC[13]); // @[bht.scala 94:27]
  wire  bhtWAddr_hash5 = io_takenPC[7] ^ (io_takenPC[13] ^ io_takenPC[14]); // @[bht.scala 95:27]
  wire  bhtWAddr_hash6 = io_takenPC[8] ^ _bhtWAddr_hash1_T_2; // @[bht.scala 96:27]
  wire [6:0] bhtWAddr = {bhtWAddr_hash6,bhtWAddr_hash5,bhtWAddr_hash4,bhtWAddr_hash3,bhtWAddr_hash2,bhtWAddr_hash1,
    bhtWAddr_hash0}; // @[bht.scala 97:58]
  wire [6:0] pht1WAddr = bhtWAddr ^ ghr; // @[bht.scala 102:26]
  wire [6:0] _GEN_897 = 7'h1 == bhtWAddr ? bht_1 : bht_0; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_898 = 7'h2 == bhtWAddr ? bht_2 : _GEN_897; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_899 = 7'h3 == bhtWAddr ? bht_3 : _GEN_898; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_900 = 7'h4 == bhtWAddr ? bht_4 : _GEN_899; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_901 = 7'h5 == bhtWAddr ? bht_5 : _GEN_900; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_902 = 7'h6 == bhtWAddr ? bht_6 : _GEN_901; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_903 = 7'h7 == bhtWAddr ? bht_7 : _GEN_902; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_904 = 7'h8 == bhtWAddr ? bht_8 : _GEN_903; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_905 = 7'h9 == bhtWAddr ? bht_9 : _GEN_904; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_906 = 7'ha == bhtWAddr ? bht_10 : _GEN_905; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_907 = 7'hb == bhtWAddr ? bht_11 : _GEN_906; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_908 = 7'hc == bhtWAddr ? bht_12 : _GEN_907; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_909 = 7'hd == bhtWAddr ? bht_13 : _GEN_908; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_910 = 7'he == bhtWAddr ? bht_14 : _GEN_909; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_911 = 7'hf == bhtWAddr ? bht_15 : _GEN_910; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_912 = 7'h10 == bhtWAddr ? bht_16 : _GEN_911; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_913 = 7'h11 == bhtWAddr ? bht_17 : _GEN_912; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_914 = 7'h12 == bhtWAddr ? bht_18 : _GEN_913; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_915 = 7'h13 == bhtWAddr ? bht_19 : _GEN_914; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_916 = 7'h14 == bhtWAddr ? bht_20 : _GEN_915; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_917 = 7'h15 == bhtWAddr ? bht_21 : _GEN_916; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_918 = 7'h16 == bhtWAddr ? bht_22 : _GEN_917; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_919 = 7'h17 == bhtWAddr ? bht_23 : _GEN_918; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_920 = 7'h18 == bhtWAddr ? bht_24 : _GEN_919; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_921 = 7'h19 == bhtWAddr ? bht_25 : _GEN_920; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_922 = 7'h1a == bhtWAddr ? bht_26 : _GEN_921; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_923 = 7'h1b == bhtWAddr ? bht_27 : _GEN_922; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_924 = 7'h1c == bhtWAddr ? bht_28 : _GEN_923; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_925 = 7'h1d == bhtWAddr ? bht_29 : _GEN_924; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_926 = 7'h1e == bhtWAddr ? bht_30 : _GEN_925; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_927 = 7'h1f == bhtWAddr ? bht_31 : _GEN_926; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_928 = 7'h20 == bhtWAddr ? bht_32 : _GEN_927; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_929 = 7'h21 == bhtWAddr ? bht_33 : _GEN_928; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_930 = 7'h22 == bhtWAddr ? bht_34 : _GEN_929; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_931 = 7'h23 == bhtWAddr ? bht_35 : _GEN_930; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_932 = 7'h24 == bhtWAddr ? bht_36 : _GEN_931; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_933 = 7'h25 == bhtWAddr ? bht_37 : _GEN_932; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_934 = 7'h26 == bhtWAddr ? bht_38 : _GEN_933; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_935 = 7'h27 == bhtWAddr ? bht_39 : _GEN_934; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_936 = 7'h28 == bhtWAddr ? bht_40 : _GEN_935; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_937 = 7'h29 == bhtWAddr ? bht_41 : _GEN_936; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_938 = 7'h2a == bhtWAddr ? bht_42 : _GEN_937; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_939 = 7'h2b == bhtWAddr ? bht_43 : _GEN_938; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_940 = 7'h2c == bhtWAddr ? bht_44 : _GEN_939; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_941 = 7'h2d == bhtWAddr ? bht_45 : _GEN_940; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_942 = 7'h2e == bhtWAddr ? bht_46 : _GEN_941; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_943 = 7'h2f == bhtWAddr ? bht_47 : _GEN_942; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_944 = 7'h30 == bhtWAddr ? bht_48 : _GEN_943; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_945 = 7'h31 == bhtWAddr ? bht_49 : _GEN_944; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_946 = 7'h32 == bhtWAddr ? bht_50 : _GEN_945; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_947 = 7'h33 == bhtWAddr ? bht_51 : _GEN_946; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_948 = 7'h34 == bhtWAddr ? bht_52 : _GEN_947; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_949 = 7'h35 == bhtWAddr ? bht_53 : _GEN_948; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_950 = 7'h36 == bhtWAddr ? bht_54 : _GEN_949; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_951 = 7'h37 == bhtWAddr ? bht_55 : _GEN_950; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_952 = 7'h38 == bhtWAddr ? bht_56 : _GEN_951; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_953 = 7'h39 == bhtWAddr ? bht_57 : _GEN_952; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_954 = 7'h3a == bhtWAddr ? bht_58 : _GEN_953; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_955 = 7'h3b == bhtWAddr ? bht_59 : _GEN_954; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_956 = 7'h3c == bhtWAddr ? bht_60 : _GEN_955; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_957 = 7'h3d == bhtWAddr ? bht_61 : _GEN_956; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_958 = 7'h3e == bhtWAddr ? bht_62 : _GEN_957; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_959 = 7'h3f == bhtWAddr ? bht_63 : _GEN_958; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_960 = 7'h40 == bhtWAddr ? bht_64 : _GEN_959; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_961 = 7'h41 == bhtWAddr ? bht_65 : _GEN_960; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_962 = 7'h42 == bhtWAddr ? bht_66 : _GEN_961; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_963 = 7'h43 == bhtWAddr ? bht_67 : _GEN_962; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_964 = 7'h44 == bhtWAddr ? bht_68 : _GEN_963; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_965 = 7'h45 == bhtWAddr ? bht_69 : _GEN_964; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_966 = 7'h46 == bhtWAddr ? bht_70 : _GEN_965; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_967 = 7'h47 == bhtWAddr ? bht_71 : _GEN_966; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_968 = 7'h48 == bhtWAddr ? bht_72 : _GEN_967; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_969 = 7'h49 == bhtWAddr ? bht_73 : _GEN_968; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_970 = 7'h4a == bhtWAddr ? bht_74 : _GEN_969; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_971 = 7'h4b == bhtWAddr ? bht_75 : _GEN_970; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_972 = 7'h4c == bhtWAddr ? bht_76 : _GEN_971; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_973 = 7'h4d == bhtWAddr ? bht_77 : _GEN_972; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_974 = 7'h4e == bhtWAddr ? bht_78 : _GEN_973; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_975 = 7'h4f == bhtWAddr ? bht_79 : _GEN_974; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_976 = 7'h50 == bhtWAddr ? bht_80 : _GEN_975; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_977 = 7'h51 == bhtWAddr ? bht_81 : _GEN_976; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_978 = 7'h52 == bhtWAddr ? bht_82 : _GEN_977; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_979 = 7'h53 == bhtWAddr ? bht_83 : _GEN_978; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_980 = 7'h54 == bhtWAddr ? bht_84 : _GEN_979; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_981 = 7'h55 == bhtWAddr ? bht_85 : _GEN_980; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_982 = 7'h56 == bhtWAddr ? bht_86 : _GEN_981; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_983 = 7'h57 == bhtWAddr ? bht_87 : _GEN_982; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_984 = 7'h58 == bhtWAddr ? bht_88 : _GEN_983; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_985 = 7'h59 == bhtWAddr ? bht_89 : _GEN_984; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_986 = 7'h5a == bhtWAddr ? bht_90 : _GEN_985; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_987 = 7'h5b == bhtWAddr ? bht_91 : _GEN_986; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_988 = 7'h5c == bhtWAddr ? bht_92 : _GEN_987; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_989 = 7'h5d == bhtWAddr ? bht_93 : _GEN_988; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_990 = 7'h5e == bhtWAddr ? bht_94 : _GEN_989; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_991 = 7'h5f == bhtWAddr ? bht_95 : _GEN_990; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_992 = 7'h60 == bhtWAddr ? bht_96 : _GEN_991; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_993 = 7'h61 == bhtWAddr ? bht_97 : _GEN_992; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_994 = 7'h62 == bhtWAddr ? bht_98 : _GEN_993; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_995 = 7'h63 == bhtWAddr ? bht_99 : _GEN_994; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_996 = 7'h64 == bhtWAddr ? bht_100 : _GEN_995; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_997 = 7'h65 == bhtWAddr ? bht_101 : _GEN_996; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_998 = 7'h66 == bhtWAddr ? bht_102 : _GEN_997; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_999 = 7'h67 == bhtWAddr ? bht_103 : _GEN_998; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_1000 = 7'h68 == bhtWAddr ? bht_104 : _GEN_999; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_1001 = 7'h69 == bhtWAddr ? bht_105 : _GEN_1000; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_1002 = 7'h6a == bhtWAddr ? bht_106 : _GEN_1001; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_1003 = 7'h6b == bhtWAddr ? bht_107 : _GEN_1002; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_1004 = 7'h6c == bhtWAddr ? bht_108 : _GEN_1003; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_1005 = 7'h6d == bhtWAddr ? bht_109 : _GEN_1004; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_1006 = 7'h6e == bhtWAddr ? bht_110 : _GEN_1005; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_1007 = 7'h6f == bhtWAddr ? bht_111 : _GEN_1006; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_1008 = 7'h70 == bhtWAddr ? bht_112 : _GEN_1007; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_1009 = 7'h71 == bhtWAddr ? bht_113 : _GEN_1008; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_1010 = 7'h72 == bhtWAddr ? bht_114 : _GEN_1009; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_1011 = 7'h73 == bhtWAddr ? bht_115 : _GEN_1010; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_1012 = 7'h74 == bhtWAddr ? bht_116 : _GEN_1011; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_1013 = 7'h75 == bhtWAddr ? bht_117 : _GEN_1012; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_1014 = 7'h76 == bhtWAddr ? bht_118 : _GEN_1013; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_1015 = 7'h77 == bhtWAddr ? bht_119 : _GEN_1014; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_1016 = 7'h78 == bhtWAddr ? bht_120 : _GEN_1015; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_1017 = 7'h79 == bhtWAddr ? bht_121 : _GEN_1016; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_1018 = 7'h7a == bhtWAddr ? bht_122 : _GEN_1017; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_1019 = 7'h7b == bhtWAddr ? bht_123 : _GEN_1018; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_1020 = 7'h7c == bhtWAddr ? bht_124 : _GEN_1019; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_1021 = 7'h7d == bhtWAddr ? bht_125 : _GEN_1020; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_1022 = 7'h7e == bhtWAddr ? bht_126 : _GEN_1021; // @[bht.scala 102:{26,26}]
  wire [6:0] _GEN_1023 = 7'h7f == bhtWAddr ? bht_127 : _GEN_1022; // @[bht.scala 102:{26,26}]
  wire [6:0] pht2WAddr = bhtWAddr ^ _GEN_1023; // @[bht.scala 102:26]
  wire [1:0] _GEN_1025 = 7'h1 == pht1WAddr ? pht_1_1 : pht_1_0; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1026 = 7'h2 == pht1WAddr ? pht_1_2 : _GEN_1025; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1027 = 7'h3 == pht1WAddr ? pht_1_3 : _GEN_1026; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1028 = 7'h4 == pht1WAddr ? pht_1_4 : _GEN_1027; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1029 = 7'h5 == pht1WAddr ? pht_1_5 : _GEN_1028; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1030 = 7'h6 == pht1WAddr ? pht_1_6 : _GEN_1029; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1031 = 7'h7 == pht1WAddr ? pht_1_7 : _GEN_1030; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1032 = 7'h8 == pht1WAddr ? pht_1_8 : _GEN_1031; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1033 = 7'h9 == pht1WAddr ? pht_1_9 : _GEN_1032; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1034 = 7'ha == pht1WAddr ? pht_1_10 : _GEN_1033; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1035 = 7'hb == pht1WAddr ? pht_1_11 : _GEN_1034; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1036 = 7'hc == pht1WAddr ? pht_1_12 : _GEN_1035; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1037 = 7'hd == pht1WAddr ? pht_1_13 : _GEN_1036; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1038 = 7'he == pht1WAddr ? pht_1_14 : _GEN_1037; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1039 = 7'hf == pht1WAddr ? pht_1_15 : _GEN_1038; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1040 = 7'h10 == pht1WAddr ? pht_1_16 : _GEN_1039; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1041 = 7'h11 == pht1WAddr ? pht_1_17 : _GEN_1040; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1042 = 7'h12 == pht1WAddr ? pht_1_18 : _GEN_1041; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1043 = 7'h13 == pht1WAddr ? pht_1_19 : _GEN_1042; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1044 = 7'h14 == pht1WAddr ? pht_1_20 : _GEN_1043; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1045 = 7'h15 == pht1WAddr ? pht_1_21 : _GEN_1044; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1046 = 7'h16 == pht1WAddr ? pht_1_22 : _GEN_1045; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1047 = 7'h17 == pht1WAddr ? pht_1_23 : _GEN_1046; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1048 = 7'h18 == pht1WAddr ? pht_1_24 : _GEN_1047; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1049 = 7'h19 == pht1WAddr ? pht_1_25 : _GEN_1048; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1050 = 7'h1a == pht1WAddr ? pht_1_26 : _GEN_1049; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1051 = 7'h1b == pht1WAddr ? pht_1_27 : _GEN_1050; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1052 = 7'h1c == pht1WAddr ? pht_1_28 : _GEN_1051; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1053 = 7'h1d == pht1WAddr ? pht_1_29 : _GEN_1052; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1054 = 7'h1e == pht1WAddr ? pht_1_30 : _GEN_1053; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1055 = 7'h1f == pht1WAddr ? pht_1_31 : _GEN_1054; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1056 = 7'h20 == pht1WAddr ? pht_1_32 : _GEN_1055; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1057 = 7'h21 == pht1WAddr ? pht_1_33 : _GEN_1056; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1058 = 7'h22 == pht1WAddr ? pht_1_34 : _GEN_1057; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1059 = 7'h23 == pht1WAddr ? pht_1_35 : _GEN_1058; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1060 = 7'h24 == pht1WAddr ? pht_1_36 : _GEN_1059; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1061 = 7'h25 == pht1WAddr ? pht_1_37 : _GEN_1060; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1062 = 7'h26 == pht1WAddr ? pht_1_38 : _GEN_1061; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1063 = 7'h27 == pht1WAddr ? pht_1_39 : _GEN_1062; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1064 = 7'h28 == pht1WAddr ? pht_1_40 : _GEN_1063; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1065 = 7'h29 == pht1WAddr ? pht_1_41 : _GEN_1064; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1066 = 7'h2a == pht1WAddr ? pht_1_42 : _GEN_1065; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1067 = 7'h2b == pht1WAddr ? pht_1_43 : _GEN_1066; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1068 = 7'h2c == pht1WAddr ? pht_1_44 : _GEN_1067; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1069 = 7'h2d == pht1WAddr ? pht_1_45 : _GEN_1068; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1070 = 7'h2e == pht1WAddr ? pht_1_46 : _GEN_1069; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1071 = 7'h2f == pht1WAddr ? pht_1_47 : _GEN_1070; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1072 = 7'h30 == pht1WAddr ? pht_1_48 : _GEN_1071; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1073 = 7'h31 == pht1WAddr ? pht_1_49 : _GEN_1072; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1074 = 7'h32 == pht1WAddr ? pht_1_50 : _GEN_1073; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1075 = 7'h33 == pht1WAddr ? pht_1_51 : _GEN_1074; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1076 = 7'h34 == pht1WAddr ? pht_1_52 : _GEN_1075; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1077 = 7'h35 == pht1WAddr ? pht_1_53 : _GEN_1076; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1078 = 7'h36 == pht1WAddr ? pht_1_54 : _GEN_1077; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1079 = 7'h37 == pht1WAddr ? pht_1_55 : _GEN_1078; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1080 = 7'h38 == pht1WAddr ? pht_1_56 : _GEN_1079; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1081 = 7'h39 == pht1WAddr ? pht_1_57 : _GEN_1080; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1082 = 7'h3a == pht1WAddr ? pht_1_58 : _GEN_1081; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1083 = 7'h3b == pht1WAddr ? pht_1_59 : _GEN_1082; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1084 = 7'h3c == pht1WAddr ? pht_1_60 : _GEN_1083; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1085 = 7'h3d == pht1WAddr ? pht_1_61 : _GEN_1084; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1086 = 7'h3e == pht1WAddr ? pht_1_62 : _GEN_1085; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1087 = 7'h3f == pht1WAddr ? pht_1_63 : _GEN_1086; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1088 = 7'h40 == pht1WAddr ? pht_1_64 : _GEN_1087; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1089 = 7'h41 == pht1WAddr ? pht_1_65 : _GEN_1088; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1090 = 7'h42 == pht1WAddr ? pht_1_66 : _GEN_1089; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1091 = 7'h43 == pht1WAddr ? pht_1_67 : _GEN_1090; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1092 = 7'h44 == pht1WAddr ? pht_1_68 : _GEN_1091; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1093 = 7'h45 == pht1WAddr ? pht_1_69 : _GEN_1092; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1094 = 7'h46 == pht1WAddr ? pht_1_70 : _GEN_1093; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1095 = 7'h47 == pht1WAddr ? pht_1_71 : _GEN_1094; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1096 = 7'h48 == pht1WAddr ? pht_1_72 : _GEN_1095; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1097 = 7'h49 == pht1WAddr ? pht_1_73 : _GEN_1096; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1098 = 7'h4a == pht1WAddr ? pht_1_74 : _GEN_1097; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1099 = 7'h4b == pht1WAddr ? pht_1_75 : _GEN_1098; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1100 = 7'h4c == pht1WAddr ? pht_1_76 : _GEN_1099; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1101 = 7'h4d == pht1WAddr ? pht_1_77 : _GEN_1100; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1102 = 7'h4e == pht1WAddr ? pht_1_78 : _GEN_1101; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1103 = 7'h4f == pht1WAddr ? pht_1_79 : _GEN_1102; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1104 = 7'h50 == pht1WAddr ? pht_1_80 : _GEN_1103; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1105 = 7'h51 == pht1WAddr ? pht_1_81 : _GEN_1104; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1106 = 7'h52 == pht1WAddr ? pht_1_82 : _GEN_1105; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1107 = 7'h53 == pht1WAddr ? pht_1_83 : _GEN_1106; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1108 = 7'h54 == pht1WAddr ? pht_1_84 : _GEN_1107; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1109 = 7'h55 == pht1WAddr ? pht_1_85 : _GEN_1108; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1110 = 7'h56 == pht1WAddr ? pht_1_86 : _GEN_1109; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1111 = 7'h57 == pht1WAddr ? pht_1_87 : _GEN_1110; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1112 = 7'h58 == pht1WAddr ? pht_1_88 : _GEN_1111; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1113 = 7'h59 == pht1WAddr ? pht_1_89 : _GEN_1112; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1114 = 7'h5a == pht1WAddr ? pht_1_90 : _GEN_1113; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1115 = 7'h5b == pht1WAddr ? pht_1_91 : _GEN_1114; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1116 = 7'h5c == pht1WAddr ? pht_1_92 : _GEN_1115; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1117 = 7'h5d == pht1WAddr ? pht_1_93 : _GEN_1116; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1118 = 7'h5e == pht1WAddr ? pht_1_94 : _GEN_1117; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1119 = 7'h5f == pht1WAddr ? pht_1_95 : _GEN_1118; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1120 = 7'h60 == pht1WAddr ? pht_1_96 : _GEN_1119; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1121 = 7'h61 == pht1WAddr ? pht_1_97 : _GEN_1120; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1122 = 7'h62 == pht1WAddr ? pht_1_98 : _GEN_1121; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1123 = 7'h63 == pht1WAddr ? pht_1_99 : _GEN_1122; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1124 = 7'h64 == pht1WAddr ? pht_1_100 : _GEN_1123; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1125 = 7'h65 == pht1WAddr ? pht_1_101 : _GEN_1124; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1126 = 7'h66 == pht1WAddr ? pht_1_102 : _GEN_1125; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1127 = 7'h67 == pht1WAddr ? pht_1_103 : _GEN_1126; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1128 = 7'h68 == pht1WAddr ? pht_1_104 : _GEN_1127; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1129 = 7'h69 == pht1WAddr ? pht_1_105 : _GEN_1128; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1130 = 7'h6a == pht1WAddr ? pht_1_106 : _GEN_1129; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1131 = 7'h6b == pht1WAddr ? pht_1_107 : _GEN_1130; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1132 = 7'h6c == pht1WAddr ? pht_1_108 : _GEN_1131; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1133 = 7'h6d == pht1WAddr ? pht_1_109 : _GEN_1132; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1134 = 7'h6e == pht1WAddr ? pht_1_110 : _GEN_1133; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1135 = 7'h6f == pht1WAddr ? pht_1_111 : _GEN_1134; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1136 = 7'h70 == pht1WAddr ? pht_1_112 : _GEN_1135; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1137 = 7'h71 == pht1WAddr ? pht_1_113 : _GEN_1136; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1138 = 7'h72 == pht1WAddr ? pht_1_114 : _GEN_1137; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1139 = 7'h73 == pht1WAddr ? pht_1_115 : _GEN_1138; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1140 = 7'h74 == pht1WAddr ? pht_1_116 : _GEN_1139; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1141 = 7'h75 == pht1WAddr ? pht_1_117 : _GEN_1140; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1142 = 7'h76 == pht1WAddr ? pht_1_118 : _GEN_1141; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1143 = 7'h77 == pht1WAddr ? pht_1_119 : _GEN_1142; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1144 = 7'h78 == pht1WAddr ? pht_1_120 : _GEN_1143; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1145 = 7'h79 == pht1WAddr ? pht_1_121 : _GEN_1144; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1146 = 7'h7a == pht1WAddr ? pht_1_122 : _GEN_1145; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1147 = 7'h7b == pht1WAddr ? pht_1_123 : _GEN_1146; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1148 = 7'h7c == pht1WAddr ? pht_1_124 : _GEN_1147; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1149 = 7'h7d == pht1WAddr ? pht_1_125 : _GEN_1148; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1150 = 7'h7e == pht1WAddr ? pht_1_126 : _GEN_1149; // @[bht.scala 156:{26,26}]
  wire [1:0] _GEN_1151 = 7'h7f == pht1WAddr ? pht_1_127 : _GEN_1150; // @[bht.scala 156:{26,26}]
  wire  p1Suc = _GEN_1151[1] == io_exTakenPre; // @[bht.scala 156:39]
  wire [1:0] _GEN_1153 = 7'h1 == pht2WAddr ? pht_2_1 : pht_2_0; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1154 = 7'h2 == pht2WAddr ? pht_2_2 : _GEN_1153; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1155 = 7'h3 == pht2WAddr ? pht_2_3 : _GEN_1154; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1156 = 7'h4 == pht2WAddr ? pht_2_4 : _GEN_1155; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1157 = 7'h5 == pht2WAddr ? pht_2_5 : _GEN_1156; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1158 = 7'h6 == pht2WAddr ? pht_2_6 : _GEN_1157; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1159 = 7'h7 == pht2WAddr ? pht_2_7 : _GEN_1158; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1160 = 7'h8 == pht2WAddr ? pht_2_8 : _GEN_1159; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1161 = 7'h9 == pht2WAddr ? pht_2_9 : _GEN_1160; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1162 = 7'ha == pht2WAddr ? pht_2_10 : _GEN_1161; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1163 = 7'hb == pht2WAddr ? pht_2_11 : _GEN_1162; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1164 = 7'hc == pht2WAddr ? pht_2_12 : _GEN_1163; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1165 = 7'hd == pht2WAddr ? pht_2_13 : _GEN_1164; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1166 = 7'he == pht2WAddr ? pht_2_14 : _GEN_1165; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1167 = 7'hf == pht2WAddr ? pht_2_15 : _GEN_1166; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1168 = 7'h10 == pht2WAddr ? pht_2_16 : _GEN_1167; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1169 = 7'h11 == pht2WAddr ? pht_2_17 : _GEN_1168; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1170 = 7'h12 == pht2WAddr ? pht_2_18 : _GEN_1169; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1171 = 7'h13 == pht2WAddr ? pht_2_19 : _GEN_1170; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1172 = 7'h14 == pht2WAddr ? pht_2_20 : _GEN_1171; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1173 = 7'h15 == pht2WAddr ? pht_2_21 : _GEN_1172; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1174 = 7'h16 == pht2WAddr ? pht_2_22 : _GEN_1173; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1175 = 7'h17 == pht2WAddr ? pht_2_23 : _GEN_1174; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1176 = 7'h18 == pht2WAddr ? pht_2_24 : _GEN_1175; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1177 = 7'h19 == pht2WAddr ? pht_2_25 : _GEN_1176; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1178 = 7'h1a == pht2WAddr ? pht_2_26 : _GEN_1177; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1179 = 7'h1b == pht2WAddr ? pht_2_27 : _GEN_1178; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1180 = 7'h1c == pht2WAddr ? pht_2_28 : _GEN_1179; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1181 = 7'h1d == pht2WAddr ? pht_2_29 : _GEN_1180; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1182 = 7'h1e == pht2WAddr ? pht_2_30 : _GEN_1181; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1183 = 7'h1f == pht2WAddr ? pht_2_31 : _GEN_1182; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1184 = 7'h20 == pht2WAddr ? pht_2_32 : _GEN_1183; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1185 = 7'h21 == pht2WAddr ? pht_2_33 : _GEN_1184; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1186 = 7'h22 == pht2WAddr ? pht_2_34 : _GEN_1185; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1187 = 7'h23 == pht2WAddr ? pht_2_35 : _GEN_1186; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1188 = 7'h24 == pht2WAddr ? pht_2_36 : _GEN_1187; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1189 = 7'h25 == pht2WAddr ? pht_2_37 : _GEN_1188; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1190 = 7'h26 == pht2WAddr ? pht_2_38 : _GEN_1189; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1191 = 7'h27 == pht2WAddr ? pht_2_39 : _GEN_1190; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1192 = 7'h28 == pht2WAddr ? pht_2_40 : _GEN_1191; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1193 = 7'h29 == pht2WAddr ? pht_2_41 : _GEN_1192; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1194 = 7'h2a == pht2WAddr ? pht_2_42 : _GEN_1193; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1195 = 7'h2b == pht2WAddr ? pht_2_43 : _GEN_1194; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1196 = 7'h2c == pht2WAddr ? pht_2_44 : _GEN_1195; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1197 = 7'h2d == pht2WAddr ? pht_2_45 : _GEN_1196; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1198 = 7'h2e == pht2WAddr ? pht_2_46 : _GEN_1197; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1199 = 7'h2f == pht2WAddr ? pht_2_47 : _GEN_1198; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1200 = 7'h30 == pht2WAddr ? pht_2_48 : _GEN_1199; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1201 = 7'h31 == pht2WAddr ? pht_2_49 : _GEN_1200; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1202 = 7'h32 == pht2WAddr ? pht_2_50 : _GEN_1201; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1203 = 7'h33 == pht2WAddr ? pht_2_51 : _GEN_1202; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1204 = 7'h34 == pht2WAddr ? pht_2_52 : _GEN_1203; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1205 = 7'h35 == pht2WAddr ? pht_2_53 : _GEN_1204; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1206 = 7'h36 == pht2WAddr ? pht_2_54 : _GEN_1205; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1207 = 7'h37 == pht2WAddr ? pht_2_55 : _GEN_1206; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1208 = 7'h38 == pht2WAddr ? pht_2_56 : _GEN_1207; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1209 = 7'h39 == pht2WAddr ? pht_2_57 : _GEN_1208; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1210 = 7'h3a == pht2WAddr ? pht_2_58 : _GEN_1209; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1211 = 7'h3b == pht2WAddr ? pht_2_59 : _GEN_1210; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1212 = 7'h3c == pht2WAddr ? pht_2_60 : _GEN_1211; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1213 = 7'h3d == pht2WAddr ? pht_2_61 : _GEN_1212; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1214 = 7'h3e == pht2WAddr ? pht_2_62 : _GEN_1213; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1215 = 7'h3f == pht2WAddr ? pht_2_63 : _GEN_1214; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1216 = 7'h40 == pht2WAddr ? pht_2_64 : _GEN_1215; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1217 = 7'h41 == pht2WAddr ? pht_2_65 : _GEN_1216; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1218 = 7'h42 == pht2WAddr ? pht_2_66 : _GEN_1217; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1219 = 7'h43 == pht2WAddr ? pht_2_67 : _GEN_1218; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1220 = 7'h44 == pht2WAddr ? pht_2_68 : _GEN_1219; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1221 = 7'h45 == pht2WAddr ? pht_2_69 : _GEN_1220; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1222 = 7'h46 == pht2WAddr ? pht_2_70 : _GEN_1221; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1223 = 7'h47 == pht2WAddr ? pht_2_71 : _GEN_1222; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1224 = 7'h48 == pht2WAddr ? pht_2_72 : _GEN_1223; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1225 = 7'h49 == pht2WAddr ? pht_2_73 : _GEN_1224; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1226 = 7'h4a == pht2WAddr ? pht_2_74 : _GEN_1225; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1227 = 7'h4b == pht2WAddr ? pht_2_75 : _GEN_1226; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1228 = 7'h4c == pht2WAddr ? pht_2_76 : _GEN_1227; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1229 = 7'h4d == pht2WAddr ? pht_2_77 : _GEN_1228; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1230 = 7'h4e == pht2WAddr ? pht_2_78 : _GEN_1229; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1231 = 7'h4f == pht2WAddr ? pht_2_79 : _GEN_1230; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1232 = 7'h50 == pht2WAddr ? pht_2_80 : _GEN_1231; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1233 = 7'h51 == pht2WAddr ? pht_2_81 : _GEN_1232; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1234 = 7'h52 == pht2WAddr ? pht_2_82 : _GEN_1233; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1235 = 7'h53 == pht2WAddr ? pht_2_83 : _GEN_1234; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1236 = 7'h54 == pht2WAddr ? pht_2_84 : _GEN_1235; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1237 = 7'h55 == pht2WAddr ? pht_2_85 : _GEN_1236; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1238 = 7'h56 == pht2WAddr ? pht_2_86 : _GEN_1237; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1239 = 7'h57 == pht2WAddr ? pht_2_87 : _GEN_1238; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1240 = 7'h58 == pht2WAddr ? pht_2_88 : _GEN_1239; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1241 = 7'h59 == pht2WAddr ? pht_2_89 : _GEN_1240; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1242 = 7'h5a == pht2WAddr ? pht_2_90 : _GEN_1241; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1243 = 7'h5b == pht2WAddr ? pht_2_91 : _GEN_1242; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1244 = 7'h5c == pht2WAddr ? pht_2_92 : _GEN_1243; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1245 = 7'h5d == pht2WAddr ? pht_2_93 : _GEN_1244; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1246 = 7'h5e == pht2WAddr ? pht_2_94 : _GEN_1245; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1247 = 7'h5f == pht2WAddr ? pht_2_95 : _GEN_1246; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1248 = 7'h60 == pht2WAddr ? pht_2_96 : _GEN_1247; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1249 = 7'h61 == pht2WAddr ? pht_2_97 : _GEN_1248; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1250 = 7'h62 == pht2WAddr ? pht_2_98 : _GEN_1249; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1251 = 7'h63 == pht2WAddr ? pht_2_99 : _GEN_1250; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1252 = 7'h64 == pht2WAddr ? pht_2_100 : _GEN_1251; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1253 = 7'h65 == pht2WAddr ? pht_2_101 : _GEN_1252; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1254 = 7'h66 == pht2WAddr ? pht_2_102 : _GEN_1253; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1255 = 7'h67 == pht2WAddr ? pht_2_103 : _GEN_1254; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1256 = 7'h68 == pht2WAddr ? pht_2_104 : _GEN_1255; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1257 = 7'h69 == pht2WAddr ? pht_2_105 : _GEN_1256; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1258 = 7'h6a == pht2WAddr ? pht_2_106 : _GEN_1257; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1259 = 7'h6b == pht2WAddr ? pht_2_107 : _GEN_1258; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1260 = 7'h6c == pht2WAddr ? pht_2_108 : _GEN_1259; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1261 = 7'h6d == pht2WAddr ? pht_2_109 : _GEN_1260; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1262 = 7'h6e == pht2WAddr ? pht_2_110 : _GEN_1261; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1263 = 7'h6f == pht2WAddr ? pht_2_111 : _GEN_1262; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1264 = 7'h70 == pht2WAddr ? pht_2_112 : _GEN_1263; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1265 = 7'h71 == pht2WAddr ? pht_2_113 : _GEN_1264; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1266 = 7'h72 == pht2WAddr ? pht_2_114 : _GEN_1265; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1267 = 7'h73 == pht2WAddr ? pht_2_115 : _GEN_1266; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1268 = 7'h74 == pht2WAddr ? pht_2_116 : _GEN_1267; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1269 = 7'h75 == pht2WAddr ? pht_2_117 : _GEN_1268; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1270 = 7'h76 == pht2WAddr ? pht_2_118 : _GEN_1269; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1271 = 7'h77 == pht2WAddr ? pht_2_119 : _GEN_1270; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1272 = 7'h78 == pht2WAddr ? pht_2_120 : _GEN_1271; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1273 = 7'h79 == pht2WAddr ? pht_2_121 : _GEN_1272; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1274 = 7'h7a == pht2WAddr ? pht_2_122 : _GEN_1273; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1275 = 7'h7b == pht2WAddr ? pht_2_123 : _GEN_1274; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1276 = 7'h7c == pht2WAddr ? pht_2_124 : _GEN_1275; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1277 = 7'h7d == pht2WAddr ? pht_2_125 : _GEN_1276; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1278 = 7'h7e == pht2WAddr ? pht_2_126 : _GEN_1277; // @[bht.scala 157:{26,26}]
  wire [1:0] _GEN_1279 = 7'h7f == pht2WAddr ? pht_2_127 : _GEN_1278; // @[bht.scala 157:{26,26}]
  wire  p2Suc = _GEN_1279[1] == io_exTakenPre; // @[bht.scala 157:39]
  wire [1:0] pht0Choice = {p1Suc,p2Suc}; // @[bht.scala 158:28]
  wire  _T = io_fire & io_takenValid; // @[bht.scala 161:18]
  wire  _pht_0_T = pht0Choice == 2'h1; // @[bht.scala 163:35]
  wire  _pht_0_T_3 = pht0Choice == 2'h2; // @[bht.scala 165:38]
  wire  _pht_0_T_4 = pht0Choice == 2'h2 ? 1'h0 : 1'h1; // @[bht.scala 165:26]
  wire [1:0] _pht_0_T_5 = _pht_0_T ? 2'h2 : {{1'd0}, _pht_0_T_4}; // @[bht.scala 164:23]
  wire [1:0] _pht_0_T_8 = _pht_0_T ? 2'h3 : 2'h2; // @[bht.scala 167:26]
  wire [1:0] _pht_0_T_9 = _pht_0_T_3 ? 2'h1 : _pht_0_T_8; // @[bht.scala 166:23]
  wire [1:0] _pht_0_T_11 = _pht_0_T_3 ? 2'h2 : 2'h3; // @[bht.scala 168:23]
  wire [1:0] _GEN_1281 = 7'h1 == pht1WAddr ? pht_0_1 : pht_0_0; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1282 = 7'h2 == pht1WAddr ? pht_0_2 : _GEN_1281; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1283 = 7'h3 == pht1WAddr ? pht_0_3 : _GEN_1282; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1284 = 7'h4 == pht1WAddr ? pht_0_4 : _GEN_1283; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1285 = 7'h5 == pht1WAddr ? pht_0_5 : _GEN_1284; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1286 = 7'h6 == pht1WAddr ? pht_0_6 : _GEN_1285; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1287 = 7'h7 == pht1WAddr ? pht_0_7 : _GEN_1286; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1288 = 7'h8 == pht1WAddr ? pht_0_8 : _GEN_1287; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1289 = 7'h9 == pht1WAddr ? pht_0_9 : _GEN_1288; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1290 = 7'ha == pht1WAddr ? pht_0_10 : _GEN_1289; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1291 = 7'hb == pht1WAddr ? pht_0_11 : _GEN_1290; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1292 = 7'hc == pht1WAddr ? pht_0_12 : _GEN_1291; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1293 = 7'hd == pht1WAddr ? pht_0_13 : _GEN_1292; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1294 = 7'he == pht1WAddr ? pht_0_14 : _GEN_1293; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1295 = 7'hf == pht1WAddr ? pht_0_15 : _GEN_1294; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1296 = 7'h10 == pht1WAddr ? pht_0_16 : _GEN_1295; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1297 = 7'h11 == pht1WAddr ? pht_0_17 : _GEN_1296; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1298 = 7'h12 == pht1WAddr ? pht_0_18 : _GEN_1297; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1299 = 7'h13 == pht1WAddr ? pht_0_19 : _GEN_1298; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1300 = 7'h14 == pht1WAddr ? pht_0_20 : _GEN_1299; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1301 = 7'h15 == pht1WAddr ? pht_0_21 : _GEN_1300; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1302 = 7'h16 == pht1WAddr ? pht_0_22 : _GEN_1301; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1303 = 7'h17 == pht1WAddr ? pht_0_23 : _GEN_1302; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1304 = 7'h18 == pht1WAddr ? pht_0_24 : _GEN_1303; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1305 = 7'h19 == pht1WAddr ? pht_0_25 : _GEN_1304; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1306 = 7'h1a == pht1WAddr ? pht_0_26 : _GEN_1305; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1307 = 7'h1b == pht1WAddr ? pht_0_27 : _GEN_1306; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1308 = 7'h1c == pht1WAddr ? pht_0_28 : _GEN_1307; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1309 = 7'h1d == pht1WAddr ? pht_0_29 : _GEN_1308; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1310 = 7'h1e == pht1WAddr ? pht_0_30 : _GEN_1309; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1311 = 7'h1f == pht1WAddr ? pht_0_31 : _GEN_1310; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1312 = 7'h20 == pht1WAddr ? pht_0_32 : _GEN_1311; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1313 = 7'h21 == pht1WAddr ? pht_0_33 : _GEN_1312; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1314 = 7'h22 == pht1WAddr ? pht_0_34 : _GEN_1313; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1315 = 7'h23 == pht1WAddr ? pht_0_35 : _GEN_1314; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1316 = 7'h24 == pht1WAddr ? pht_0_36 : _GEN_1315; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1317 = 7'h25 == pht1WAddr ? pht_0_37 : _GEN_1316; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1318 = 7'h26 == pht1WAddr ? pht_0_38 : _GEN_1317; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1319 = 7'h27 == pht1WAddr ? pht_0_39 : _GEN_1318; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1320 = 7'h28 == pht1WAddr ? pht_0_40 : _GEN_1319; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1321 = 7'h29 == pht1WAddr ? pht_0_41 : _GEN_1320; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1322 = 7'h2a == pht1WAddr ? pht_0_42 : _GEN_1321; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1323 = 7'h2b == pht1WAddr ? pht_0_43 : _GEN_1322; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1324 = 7'h2c == pht1WAddr ? pht_0_44 : _GEN_1323; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1325 = 7'h2d == pht1WAddr ? pht_0_45 : _GEN_1324; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1326 = 7'h2e == pht1WAddr ? pht_0_46 : _GEN_1325; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1327 = 7'h2f == pht1WAddr ? pht_0_47 : _GEN_1326; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1328 = 7'h30 == pht1WAddr ? pht_0_48 : _GEN_1327; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1329 = 7'h31 == pht1WAddr ? pht_0_49 : _GEN_1328; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1330 = 7'h32 == pht1WAddr ? pht_0_50 : _GEN_1329; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1331 = 7'h33 == pht1WAddr ? pht_0_51 : _GEN_1330; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1332 = 7'h34 == pht1WAddr ? pht_0_52 : _GEN_1331; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1333 = 7'h35 == pht1WAddr ? pht_0_53 : _GEN_1332; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1334 = 7'h36 == pht1WAddr ? pht_0_54 : _GEN_1333; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1335 = 7'h37 == pht1WAddr ? pht_0_55 : _GEN_1334; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1336 = 7'h38 == pht1WAddr ? pht_0_56 : _GEN_1335; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1337 = 7'h39 == pht1WAddr ? pht_0_57 : _GEN_1336; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1338 = 7'h3a == pht1WAddr ? pht_0_58 : _GEN_1337; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1339 = 7'h3b == pht1WAddr ? pht_0_59 : _GEN_1338; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1340 = 7'h3c == pht1WAddr ? pht_0_60 : _GEN_1339; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1341 = 7'h3d == pht1WAddr ? pht_0_61 : _GEN_1340; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1342 = 7'h3e == pht1WAddr ? pht_0_62 : _GEN_1341; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1343 = 7'h3f == pht1WAddr ? pht_0_63 : _GEN_1342; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1344 = 7'h40 == pht1WAddr ? pht_0_64 : _GEN_1343; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1345 = 7'h41 == pht1WAddr ? pht_0_65 : _GEN_1344; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1346 = 7'h42 == pht1WAddr ? pht_0_66 : _GEN_1345; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1347 = 7'h43 == pht1WAddr ? pht_0_67 : _GEN_1346; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1348 = 7'h44 == pht1WAddr ? pht_0_68 : _GEN_1347; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1349 = 7'h45 == pht1WAddr ? pht_0_69 : _GEN_1348; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1350 = 7'h46 == pht1WAddr ? pht_0_70 : _GEN_1349; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1351 = 7'h47 == pht1WAddr ? pht_0_71 : _GEN_1350; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1352 = 7'h48 == pht1WAddr ? pht_0_72 : _GEN_1351; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1353 = 7'h49 == pht1WAddr ? pht_0_73 : _GEN_1352; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1354 = 7'h4a == pht1WAddr ? pht_0_74 : _GEN_1353; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1355 = 7'h4b == pht1WAddr ? pht_0_75 : _GEN_1354; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1356 = 7'h4c == pht1WAddr ? pht_0_76 : _GEN_1355; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1357 = 7'h4d == pht1WAddr ? pht_0_77 : _GEN_1356; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1358 = 7'h4e == pht1WAddr ? pht_0_78 : _GEN_1357; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1359 = 7'h4f == pht1WAddr ? pht_0_79 : _GEN_1358; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1360 = 7'h50 == pht1WAddr ? pht_0_80 : _GEN_1359; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1361 = 7'h51 == pht1WAddr ? pht_0_81 : _GEN_1360; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1362 = 7'h52 == pht1WAddr ? pht_0_82 : _GEN_1361; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1363 = 7'h53 == pht1WAddr ? pht_0_83 : _GEN_1362; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1364 = 7'h54 == pht1WAddr ? pht_0_84 : _GEN_1363; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1365 = 7'h55 == pht1WAddr ? pht_0_85 : _GEN_1364; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1366 = 7'h56 == pht1WAddr ? pht_0_86 : _GEN_1365; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1367 = 7'h57 == pht1WAddr ? pht_0_87 : _GEN_1366; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1368 = 7'h58 == pht1WAddr ? pht_0_88 : _GEN_1367; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1369 = 7'h59 == pht1WAddr ? pht_0_89 : _GEN_1368; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1370 = 7'h5a == pht1WAddr ? pht_0_90 : _GEN_1369; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1371 = 7'h5b == pht1WAddr ? pht_0_91 : _GEN_1370; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1372 = 7'h5c == pht1WAddr ? pht_0_92 : _GEN_1371; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1373 = 7'h5d == pht1WAddr ? pht_0_93 : _GEN_1372; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1374 = 7'h5e == pht1WAddr ? pht_0_94 : _GEN_1373; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1375 = 7'h5f == pht1WAddr ? pht_0_95 : _GEN_1374; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1376 = 7'h60 == pht1WAddr ? pht_0_96 : _GEN_1375; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1377 = 7'h61 == pht1WAddr ? pht_0_97 : _GEN_1376; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1378 = 7'h62 == pht1WAddr ? pht_0_98 : _GEN_1377; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1379 = 7'h63 == pht1WAddr ? pht_0_99 : _GEN_1378; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1380 = 7'h64 == pht1WAddr ? pht_0_100 : _GEN_1379; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1381 = 7'h65 == pht1WAddr ? pht_0_101 : _GEN_1380; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1382 = 7'h66 == pht1WAddr ? pht_0_102 : _GEN_1381; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1383 = 7'h67 == pht1WAddr ? pht_0_103 : _GEN_1382; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1384 = 7'h68 == pht1WAddr ? pht_0_104 : _GEN_1383; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1385 = 7'h69 == pht1WAddr ? pht_0_105 : _GEN_1384; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1386 = 7'h6a == pht1WAddr ? pht_0_106 : _GEN_1385; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1387 = 7'h6b == pht1WAddr ? pht_0_107 : _GEN_1386; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1388 = 7'h6c == pht1WAddr ? pht_0_108 : _GEN_1387; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1389 = 7'h6d == pht1WAddr ? pht_0_109 : _GEN_1388; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1390 = 7'h6e == pht1WAddr ? pht_0_110 : _GEN_1389; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1391 = 7'h6f == pht1WAddr ? pht_0_111 : _GEN_1390; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1392 = 7'h70 == pht1WAddr ? pht_0_112 : _GEN_1391; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1393 = 7'h71 == pht1WAddr ? pht_0_113 : _GEN_1392; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1394 = 7'h72 == pht1WAddr ? pht_0_114 : _GEN_1393; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1395 = 7'h73 == pht1WAddr ? pht_0_115 : _GEN_1394; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1396 = 7'h74 == pht1WAddr ? pht_0_116 : _GEN_1395; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1397 = 7'h75 == pht1WAddr ? pht_0_117 : _GEN_1396; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1398 = 7'h76 == pht1WAddr ? pht_0_118 : _GEN_1397; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1399 = 7'h77 == pht1WAddr ? pht_0_119 : _GEN_1398; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1400 = 7'h78 == pht1WAddr ? pht_0_120 : _GEN_1399; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1401 = 7'h79 == pht1WAddr ? pht_0_121 : _GEN_1400; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1402 = 7'h7a == pht1WAddr ? pht_0_122 : _GEN_1401; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1403 = 7'h7b == pht1WAddr ? pht_0_123 : _GEN_1402; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1404 = 7'h7c == pht1WAddr ? pht_0_124 : _GEN_1403; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1405 = 7'h7d == pht1WAddr ? pht_0_125 : _GEN_1404; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1406 = 7'h7e == pht1WAddr ? pht_0_126 : _GEN_1405; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1407 = 7'h7f == pht1WAddr ? pht_0_127 : _GEN_1406; // @[Mux.scala 81:{61,61}]
  wire [1:0] _pht_0_T_13 = 2'h1 == _GEN_1407 ? _pht_0_T_5 : {{1'd0}, _pht_0_T}; // @[Mux.scala 81:58]
  wire [1:0] _pht_0_T_15 = 2'h2 == _GEN_1407 ? _pht_0_T_9 : _pht_0_T_13; // @[Mux.scala 81:58]
  wire [1:0] _pht_1_T_1 = io_takenMiss ? 2'h2 : 2'h0; // @[bht.scala 174:23]
  wire [1:0] _pht_1_T_2 = io_takenMiss ? 2'h1 : 2'h3; // @[bht.scala 175:23]
  wire [1:0] _pht_1_T_3 = io_takenMiss ? 2'h2 : 2'h3; // @[bht.scala 176:23]
  wire [1:0] _pht_1_T_5 = 2'h1 == _GEN_1151 ? _pht_1_T_1 : {{1'd0}, io_takenMiss}; // @[Mux.scala 81:58]
  wire [1:0] _pht_1_T_7 = 2'h2 == _GEN_1151 ? _pht_1_T_2 : _pht_1_T_5; // @[Mux.scala 81:58]
  wire [1:0] _pht_2_T_5 = 2'h1 == _GEN_1279 ? _pht_1_T_1 : {{1'd0}, io_takenMiss}; // @[Mux.scala 81:58]
  wire [1:0] _pht_2_T_7 = 2'h2 == _GEN_1279 ? _pht_1_T_2 : _pht_2_T_5; // @[Mux.scala 81:58]
  wire [6:0] _bht_T_1 = {_GEN_1023[5:0],io_exTakenPre}; // @[bht.scala 189:49]
  wire [6:0] _ghr_T_1 = {ghr[5:0],io_exTakenPre}; // @[bht.scala 190:33]
  wire [6:0] upIndex = io_takenPC[10:4]; // @[bht.scala 194:27]
  wire  _GEN_2433 = 7'h0 == upIndex | btbV_0; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2434 = 7'h1 == upIndex | btbV_1; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2435 = 7'h2 == upIndex | btbV_2; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2436 = 7'h3 == upIndex | btbV_3; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2437 = 7'h4 == upIndex | btbV_4; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2438 = 7'h5 == upIndex | btbV_5; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2439 = 7'h6 == upIndex | btbV_6; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2440 = 7'h7 == upIndex | btbV_7; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2441 = 7'h8 == upIndex | btbV_8; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2442 = 7'h9 == upIndex | btbV_9; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2443 = 7'ha == upIndex | btbV_10; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2444 = 7'hb == upIndex | btbV_11; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2445 = 7'hc == upIndex | btbV_12; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2446 = 7'hd == upIndex | btbV_13; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2447 = 7'he == upIndex | btbV_14; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2448 = 7'hf == upIndex | btbV_15; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2449 = 7'h10 == upIndex | btbV_16; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2450 = 7'h11 == upIndex | btbV_17; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2451 = 7'h12 == upIndex | btbV_18; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2452 = 7'h13 == upIndex | btbV_19; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2453 = 7'h14 == upIndex | btbV_20; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2454 = 7'h15 == upIndex | btbV_21; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2455 = 7'h16 == upIndex | btbV_22; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2456 = 7'h17 == upIndex | btbV_23; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2457 = 7'h18 == upIndex | btbV_24; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2458 = 7'h19 == upIndex | btbV_25; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2459 = 7'h1a == upIndex | btbV_26; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2460 = 7'h1b == upIndex | btbV_27; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2461 = 7'h1c == upIndex | btbV_28; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2462 = 7'h1d == upIndex | btbV_29; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2463 = 7'h1e == upIndex | btbV_30; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2464 = 7'h1f == upIndex | btbV_31; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2465 = 7'h20 == upIndex | btbV_32; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2466 = 7'h21 == upIndex | btbV_33; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2467 = 7'h22 == upIndex | btbV_34; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2468 = 7'h23 == upIndex | btbV_35; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2469 = 7'h24 == upIndex | btbV_36; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2470 = 7'h25 == upIndex | btbV_37; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2471 = 7'h26 == upIndex | btbV_38; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2472 = 7'h27 == upIndex | btbV_39; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2473 = 7'h28 == upIndex | btbV_40; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2474 = 7'h29 == upIndex | btbV_41; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2475 = 7'h2a == upIndex | btbV_42; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2476 = 7'h2b == upIndex | btbV_43; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2477 = 7'h2c == upIndex | btbV_44; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2478 = 7'h2d == upIndex | btbV_45; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2479 = 7'h2e == upIndex | btbV_46; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2480 = 7'h2f == upIndex | btbV_47; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2481 = 7'h30 == upIndex | btbV_48; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2482 = 7'h31 == upIndex | btbV_49; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2483 = 7'h32 == upIndex | btbV_50; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2484 = 7'h33 == upIndex | btbV_51; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2485 = 7'h34 == upIndex | btbV_52; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2486 = 7'h35 == upIndex | btbV_53; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2487 = 7'h36 == upIndex | btbV_54; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2488 = 7'h37 == upIndex | btbV_55; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2489 = 7'h38 == upIndex | btbV_56; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2490 = 7'h39 == upIndex | btbV_57; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2491 = 7'h3a == upIndex | btbV_58; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2492 = 7'h3b == upIndex | btbV_59; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2493 = 7'h3c == upIndex | btbV_60; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2494 = 7'h3d == upIndex | btbV_61; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2495 = 7'h3e == upIndex | btbV_62; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2496 = 7'h3f == upIndex | btbV_63; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2497 = 7'h40 == upIndex | btbV_64; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2498 = 7'h41 == upIndex | btbV_65; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2499 = 7'h42 == upIndex | btbV_66; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2500 = 7'h43 == upIndex | btbV_67; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2501 = 7'h44 == upIndex | btbV_68; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2502 = 7'h45 == upIndex | btbV_69; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2503 = 7'h46 == upIndex | btbV_70; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2504 = 7'h47 == upIndex | btbV_71; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2505 = 7'h48 == upIndex | btbV_72; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2506 = 7'h49 == upIndex | btbV_73; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2507 = 7'h4a == upIndex | btbV_74; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2508 = 7'h4b == upIndex | btbV_75; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2509 = 7'h4c == upIndex | btbV_76; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2510 = 7'h4d == upIndex | btbV_77; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2511 = 7'h4e == upIndex | btbV_78; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2512 = 7'h4f == upIndex | btbV_79; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2513 = 7'h50 == upIndex | btbV_80; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2514 = 7'h51 == upIndex | btbV_81; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2515 = 7'h52 == upIndex | btbV_82; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2516 = 7'h53 == upIndex | btbV_83; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2517 = 7'h54 == upIndex | btbV_84; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2518 = 7'h55 == upIndex | btbV_85; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2519 = 7'h56 == upIndex | btbV_86; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2520 = 7'h57 == upIndex | btbV_87; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2521 = 7'h58 == upIndex | btbV_88; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2522 = 7'h59 == upIndex | btbV_89; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2523 = 7'h5a == upIndex | btbV_90; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2524 = 7'h5b == upIndex | btbV_91; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2525 = 7'h5c == upIndex | btbV_92; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2526 = 7'h5d == upIndex | btbV_93; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2527 = 7'h5e == upIndex | btbV_94; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2528 = 7'h5f == upIndex | btbV_95; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2529 = 7'h60 == upIndex | btbV_96; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2530 = 7'h61 == upIndex | btbV_97; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2531 = 7'h62 == upIndex | btbV_98; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2532 = 7'h63 == upIndex | btbV_99; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2533 = 7'h64 == upIndex | btbV_100; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2534 = 7'h65 == upIndex | btbV_101; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2535 = 7'h66 == upIndex | btbV_102; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2536 = 7'h67 == upIndex | btbV_103; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2537 = 7'h68 == upIndex | btbV_104; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2538 = 7'h69 == upIndex | btbV_105; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2539 = 7'h6a == upIndex | btbV_106; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2540 = 7'h6b == upIndex | btbV_107; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2541 = 7'h6c == upIndex | btbV_108; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2542 = 7'h6d == upIndex | btbV_109; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2543 = 7'h6e == upIndex | btbV_110; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2544 = 7'h6f == upIndex | btbV_111; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2545 = 7'h70 == upIndex | btbV_112; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2546 = 7'h71 == upIndex | btbV_113; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2547 = 7'h72 == upIndex | btbV_114; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2548 = 7'h73 == upIndex | btbV_115; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2549 = 7'h74 == upIndex | btbV_116; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2550 = 7'h75 == upIndex | btbV_117; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2551 = 7'h76 == upIndex | btbV_118; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2552 = 7'h77 == upIndex | btbV_119; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2553 = 7'h78 == upIndex | btbV_120; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2554 = 7'h79 == upIndex | btbV_121; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2555 = 7'h7a == upIndex | btbV_122; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2556 = 7'h7b == upIndex | btbV_123; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2557 = 7'h7c == upIndex | btbV_124; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2558 = 7'h7d == upIndex | btbV_125; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2559 = 7'h7e == upIndex | btbV_126; // @[bht.scala 198:{19,19} 112:23]
  wire  _GEN_2560 = 7'h7f == upIndex | btbV_127; // @[bht.scala 198:{19,19} 112:23]
  assign io_takenPre = io_valid & _io_takenPre_T_4; // @[bht.scala 132:23]
  assign io_takenPrePC = _io_takenPrePC_T_4[31:0]; // @[bht.scala 137:19]
  assign io_ready = io_valid & io_bxx ? io_ready_REG : io_fire; // @[bht.scala 142:20]
  always @(posedge clock) begin
    if (reset) begin // @[bht.scala 107:22]
      ghr <= 7'h0; // @[bht.scala 107:22]
    end else if (_T) begin // @[bht.scala 188:36]
      ghr <= _ghr_T_1; // @[bht.scala 190:11]
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_0 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h0 == bhtWAddr) begin // @[bht.scala 189:21]
        bht_0 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_1 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h1 == bhtWAddr) begin // @[bht.scala 189:21]
        bht_1 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_2 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h2 == bhtWAddr) begin // @[bht.scala 189:21]
        bht_2 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_3 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h3 == bhtWAddr) begin // @[bht.scala 189:21]
        bht_3 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_4 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h4 == bhtWAddr) begin // @[bht.scala 189:21]
        bht_4 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_5 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h5 == bhtWAddr) begin // @[bht.scala 189:21]
        bht_5 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_6 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h6 == bhtWAddr) begin // @[bht.scala 189:21]
        bht_6 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_7 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h7 == bhtWAddr) begin // @[bht.scala 189:21]
        bht_7 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_8 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h8 == bhtWAddr) begin // @[bht.scala 189:21]
        bht_8 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_9 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h9 == bhtWAddr) begin // @[bht.scala 189:21]
        bht_9 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_10 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'ha == bhtWAddr) begin // @[bht.scala 189:21]
        bht_10 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_11 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'hb == bhtWAddr) begin // @[bht.scala 189:21]
        bht_11 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_12 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'hc == bhtWAddr) begin // @[bht.scala 189:21]
        bht_12 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_13 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'hd == bhtWAddr) begin // @[bht.scala 189:21]
        bht_13 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_14 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'he == bhtWAddr) begin // @[bht.scala 189:21]
        bht_14 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_15 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'hf == bhtWAddr) begin // @[bht.scala 189:21]
        bht_15 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_16 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h10 == bhtWAddr) begin // @[bht.scala 189:21]
        bht_16 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_17 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h11 == bhtWAddr) begin // @[bht.scala 189:21]
        bht_17 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_18 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h12 == bhtWAddr) begin // @[bht.scala 189:21]
        bht_18 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_19 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h13 == bhtWAddr) begin // @[bht.scala 189:21]
        bht_19 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_20 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h14 == bhtWAddr) begin // @[bht.scala 189:21]
        bht_20 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_21 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h15 == bhtWAddr) begin // @[bht.scala 189:21]
        bht_21 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_22 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h16 == bhtWAddr) begin // @[bht.scala 189:21]
        bht_22 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_23 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h17 == bhtWAddr) begin // @[bht.scala 189:21]
        bht_23 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_24 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h18 == bhtWAddr) begin // @[bht.scala 189:21]
        bht_24 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_25 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h19 == bhtWAddr) begin // @[bht.scala 189:21]
        bht_25 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_26 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h1a == bhtWAddr) begin // @[bht.scala 189:21]
        bht_26 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_27 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h1b == bhtWAddr) begin // @[bht.scala 189:21]
        bht_27 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_28 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h1c == bhtWAddr) begin // @[bht.scala 189:21]
        bht_28 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_29 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h1d == bhtWAddr) begin // @[bht.scala 189:21]
        bht_29 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_30 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h1e == bhtWAddr) begin // @[bht.scala 189:21]
        bht_30 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_31 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h1f == bhtWAddr) begin // @[bht.scala 189:21]
        bht_31 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_32 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h20 == bhtWAddr) begin // @[bht.scala 189:21]
        bht_32 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_33 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h21 == bhtWAddr) begin // @[bht.scala 189:21]
        bht_33 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_34 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h22 == bhtWAddr) begin // @[bht.scala 189:21]
        bht_34 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_35 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h23 == bhtWAddr) begin // @[bht.scala 189:21]
        bht_35 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_36 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h24 == bhtWAddr) begin // @[bht.scala 189:21]
        bht_36 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_37 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h25 == bhtWAddr) begin // @[bht.scala 189:21]
        bht_37 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_38 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h26 == bhtWAddr) begin // @[bht.scala 189:21]
        bht_38 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_39 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h27 == bhtWAddr) begin // @[bht.scala 189:21]
        bht_39 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_40 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h28 == bhtWAddr) begin // @[bht.scala 189:21]
        bht_40 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_41 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h29 == bhtWAddr) begin // @[bht.scala 189:21]
        bht_41 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_42 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h2a == bhtWAddr) begin // @[bht.scala 189:21]
        bht_42 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_43 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h2b == bhtWAddr) begin // @[bht.scala 189:21]
        bht_43 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_44 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h2c == bhtWAddr) begin // @[bht.scala 189:21]
        bht_44 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_45 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h2d == bhtWAddr) begin // @[bht.scala 189:21]
        bht_45 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_46 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h2e == bhtWAddr) begin // @[bht.scala 189:21]
        bht_46 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_47 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h2f == bhtWAddr) begin // @[bht.scala 189:21]
        bht_47 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_48 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h30 == bhtWAddr) begin // @[bht.scala 189:21]
        bht_48 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_49 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h31 == bhtWAddr) begin // @[bht.scala 189:21]
        bht_49 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_50 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h32 == bhtWAddr) begin // @[bht.scala 189:21]
        bht_50 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_51 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h33 == bhtWAddr) begin // @[bht.scala 189:21]
        bht_51 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_52 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h34 == bhtWAddr) begin // @[bht.scala 189:21]
        bht_52 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_53 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h35 == bhtWAddr) begin // @[bht.scala 189:21]
        bht_53 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_54 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h36 == bhtWAddr) begin // @[bht.scala 189:21]
        bht_54 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_55 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h37 == bhtWAddr) begin // @[bht.scala 189:21]
        bht_55 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_56 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h38 == bhtWAddr) begin // @[bht.scala 189:21]
        bht_56 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_57 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h39 == bhtWAddr) begin // @[bht.scala 189:21]
        bht_57 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_58 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h3a == bhtWAddr) begin // @[bht.scala 189:21]
        bht_58 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_59 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h3b == bhtWAddr) begin // @[bht.scala 189:21]
        bht_59 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_60 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h3c == bhtWAddr) begin // @[bht.scala 189:21]
        bht_60 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_61 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h3d == bhtWAddr) begin // @[bht.scala 189:21]
        bht_61 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_62 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h3e == bhtWAddr) begin // @[bht.scala 189:21]
        bht_62 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_63 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h3f == bhtWAddr) begin // @[bht.scala 189:21]
        bht_63 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_64 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h40 == bhtWAddr) begin // @[bht.scala 189:21]
        bht_64 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_65 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h41 == bhtWAddr) begin // @[bht.scala 189:21]
        bht_65 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_66 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h42 == bhtWAddr) begin // @[bht.scala 189:21]
        bht_66 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_67 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h43 == bhtWAddr) begin // @[bht.scala 189:21]
        bht_67 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_68 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h44 == bhtWAddr) begin // @[bht.scala 189:21]
        bht_68 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_69 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h45 == bhtWAddr) begin // @[bht.scala 189:21]
        bht_69 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_70 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h46 == bhtWAddr) begin // @[bht.scala 189:21]
        bht_70 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_71 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h47 == bhtWAddr) begin // @[bht.scala 189:21]
        bht_71 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_72 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h48 == bhtWAddr) begin // @[bht.scala 189:21]
        bht_72 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_73 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h49 == bhtWAddr) begin // @[bht.scala 189:21]
        bht_73 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_74 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h4a == bhtWAddr) begin // @[bht.scala 189:21]
        bht_74 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_75 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h4b == bhtWAddr) begin // @[bht.scala 189:21]
        bht_75 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_76 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h4c == bhtWAddr) begin // @[bht.scala 189:21]
        bht_76 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_77 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h4d == bhtWAddr) begin // @[bht.scala 189:21]
        bht_77 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_78 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h4e == bhtWAddr) begin // @[bht.scala 189:21]
        bht_78 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_79 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h4f == bhtWAddr) begin // @[bht.scala 189:21]
        bht_79 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_80 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h50 == bhtWAddr) begin // @[bht.scala 189:21]
        bht_80 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_81 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h51 == bhtWAddr) begin // @[bht.scala 189:21]
        bht_81 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_82 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h52 == bhtWAddr) begin // @[bht.scala 189:21]
        bht_82 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_83 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h53 == bhtWAddr) begin // @[bht.scala 189:21]
        bht_83 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_84 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h54 == bhtWAddr) begin // @[bht.scala 189:21]
        bht_84 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_85 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h55 == bhtWAddr) begin // @[bht.scala 189:21]
        bht_85 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_86 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h56 == bhtWAddr) begin // @[bht.scala 189:21]
        bht_86 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_87 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h57 == bhtWAddr) begin // @[bht.scala 189:21]
        bht_87 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_88 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h58 == bhtWAddr) begin // @[bht.scala 189:21]
        bht_88 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_89 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h59 == bhtWAddr) begin // @[bht.scala 189:21]
        bht_89 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_90 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h5a == bhtWAddr) begin // @[bht.scala 189:21]
        bht_90 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_91 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h5b == bhtWAddr) begin // @[bht.scala 189:21]
        bht_91 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_92 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h5c == bhtWAddr) begin // @[bht.scala 189:21]
        bht_92 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_93 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h5d == bhtWAddr) begin // @[bht.scala 189:21]
        bht_93 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_94 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h5e == bhtWAddr) begin // @[bht.scala 189:21]
        bht_94 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_95 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h5f == bhtWAddr) begin // @[bht.scala 189:21]
        bht_95 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_96 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h60 == bhtWAddr) begin // @[bht.scala 189:21]
        bht_96 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_97 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h61 == bhtWAddr) begin // @[bht.scala 189:21]
        bht_97 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_98 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h62 == bhtWAddr) begin // @[bht.scala 189:21]
        bht_98 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_99 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h63 == bhtWAddr) begin // @[bht.scala 189:21]
        bht_99 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_100 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h64 == bhtWAddr) begin // @[bht.scala 189:21]
        bht_100 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_101 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h65 == bhtWAddr) begin // @[bht.scala 189:21]
        bht_101 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_102 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h66 == bhtWAddr) begin // @[bht.scala 189:21]
        bht_102 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_103 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h67 == bhtWAddr) begin // @[bht.scala 189:21]
        bht_103 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_104 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h68 == bhtWAddr) begin // @[bht.scala 189:21]
        bht_104 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_105 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h69 == bhtWAddr) begin // @[bht.scala 189:21]
        bht_105 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_106 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h6a == bhtWAddr) begin // @[bht.scala 189:21]
        bht_106 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_107 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h6b == bhtWAddr) begin // @[bht.scala 189:21]
        bht_107 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_108 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h6c == bhtWAddr) begin // @[bht.scala 189:21]
        bht_108 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_109 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h6d == bhtWAddr) begin // @[bht.scala 189:21]
        bht_109 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_110 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h6e == bhtWAddr) begin // @[bht.scala 189:21]
        bht_110 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_111 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h6f == bhtWAddr) begin // @[bht.scala 189:21]
        bht_111 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_112 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h70 == bhtWAddr) begin // @[bht.scala 189:21]
        bht_112 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_113 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h71 == bhtWAddr) begin // @[bht.scala 189:21]
        bht_113 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_114 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h72 == bhtWAddr) begin // @[bht.scala 189:21]
        bht_114 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_115 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h73 == bhtWAddr) begin // @[bht.scala 189:21]
        bht_115 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_116 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h74 == bhtWAddr) begin // @[bht.scala 189:21]
        bht_116 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_117 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h75 == bhtWAddr) begin // @[bht.scala 189:21]
        bht_117 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_118 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h76 == bhtWAddr) begin // @[bht.scala 189:21]
        bht_118 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_119 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h77 == bhtWAddr) begin // @[bht.scala 189:21]
        bht_119 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_120 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h78 == bhtWAddr) begin // @[bht.scala 189:21]
        bht_120 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_121 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h79 == bhtWAddr) begin // @[bht.scala 189:21]
        bht_121 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_122 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h7a == bhtWAddr) begin // @[bht.scala 189:21]
        bht_122 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_123 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h7b == bhtWAddr) begin // @[bht.scala 189:21]
        bht_123 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_124 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h7c == bhtWAddr) begin // @[bht.scala 189:21]
        bht_124 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_125 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h7d == bhtWAddr) begin // @[bht.scala 189:21]
        bht_125 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_126 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h7e == bhtWAddr) begin // @[bht.scala 189:21]
        bht_126 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 108:22]
      bht_127 <= 7'h0; // @[bht.scala 108:22]
    end else if (_T) begin // @[bht.scala 188:36]
      if (7'h7f == bhtWAddr) begin // @[bht.scala 189:21]
        bht_127 <= _bht_T_1; // @[bht.scala 189:21]
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_0 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h0 == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_0 <= _pht_0_T_11;
        end else begin
          pht_0_0 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_1 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h1 == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_1 <= _pht_0_T_11;
        end else begin
          pht_0_1 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_2 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h2 == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_2 <= _pht_0_T_11;
        end else begin
          pht_0_2 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_3 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h3 == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_3 <= _pht_0_T_11;
        end else begin
          pht_0_3 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_4 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h4 == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_4 <= _pht_0_T_11;
        end else begin
          pht_0_4 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_5 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h5 == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_5 <= _pht_0_T_11;
        end else begin
          pht_0_5 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_6 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h6 == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_6 <= _pht_0_T_11;
        end else begin
          pht_0_6 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_7 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h7 == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_7 <= _pht_0_T_11;
        end else begin
          pht_0_7 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_8 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h8 == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_8 <= _pht_0_T_11;
        end else begin
          pht_0_8 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_9 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h9 == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_9 <= _pht_0_T_11;
        end else begin
          pht_0_9 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_10 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'ha == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_10 <= _pht_0_T_11;
        end else begin
          pht_0_10 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_11 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'hb == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_11 <= _pht_0_T_11;
        end else begin
          pht_0_11 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_12 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'hc == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_12 <= _pht_0_T_11;
        end else begin
          pht_0_12 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_13 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'hd == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_13 <= _pht_0_T_11;
        end else begin
          pht_0_13 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_14 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'he == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_14 <= _pht_0_T_11;
        end else begin
          pht_0_14 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_15 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'hf == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_15 <= _pht_0_T_11;
        end else begin
          pht_0_15 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_16 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h10 == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_16 <= _pht_0_T_11;
        end else begin
          pht_0_16 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_17 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h11 == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_17 <= _pht_0_T_11;
        end else begin
          pht_0_17 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_18 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h12 == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_18 <= _pht_0_T_11;
        end else begin
          pht_0_18 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_19 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h13 == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_19 <= _pht_0_T_11;
        end else begin
          pht_0_19 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_20 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h14 == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_20 <= _pht_0_T_11;
        end else begin
          pht_0_20 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_21 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h15 == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_21 <= _pht_0_T_11;
        end else begin
          pht_0_21 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_22 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h16 == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_22 <= _pht_0_T_11;
        end else begin
          pht_0_22 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_23 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h17 == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_23 <= _pht_0_T_11;
        end else begin
          pht_0_23 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_24 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h18 == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_24 <= _pht_0_T_11;
        end else begin
          pht_0_24 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_25 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h19 == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_25 <= _pht_0_T_11;
        end else begin
          pht_0_25 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_26 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h1a == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_26 <= _pht_0_T_11;
        end else begin
          pht_0_26 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_27 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h1b == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_27 <= _pht_0_T_11;
        end else begin
          pht_0_27 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_28 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h1c == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_28 <= _pht_0_T_11;
        end else begin
          pht_0_28 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_29 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h1d == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_29 <= _pht_0_T_11;
        end else begin
          pht_0_29 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_30 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h1e == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_30 <= _pht_0_T_11;
        end else begin
          pht_0_30 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_31 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h1f == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_31 <= _pht_0_T_11;
        end else begin
          pht_0_31 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_32 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h20 == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_32 <= _pht_0_T_11;
        end else begin
          pht_0_32 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_33 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h21 == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_33 <= _pht_0_T_11;
        end else begin
          pht_0_33 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_34 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h22 == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_34 <= _pht_0_T_11;
        end else begin
          pht_0_34 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_35 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h23 == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_35 <= _pht_0_T_11;
        end else begin
          pht_0_35 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_36 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h24 == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_36 <= _pht_0_T_11;
        end else begin
          pht_0_36 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_37 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h25 == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_37 <= _pht_0_T_11;
        end else begin
          pht_0_37 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_38 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h26 == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_38 <= _pht_0_T_11;
        end else begin
          pht_0_38 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_39 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h27 == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_39 <= _pht_0_T_11;
        end else begin
          pht_0_39 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_40 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h28 == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_40 <= _pht_0_T_11;
        end else begin
          pht_0_40 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_41 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h29 == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_41 <= _pht_0_T_11;
        end else begin
          pht_0_41 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_42 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h2a == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_42 <= _pht_0_T_11;
        end else begin
          pht_0_42 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_43 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h2b == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_43 <= _pht_0_T_11;
        end else begin
          pht_0_43 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_44 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h2c == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_44 <= _pht_0_T_11;
        end else begin
          pht_0_44 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_45 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h2d == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_45 <= _pht_0_T_11;
        end else begin
          pht_0_45 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_46 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h2e == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_46 <= _pht_0_T_11;
        end else begin
          pht_0_46 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_47 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h2f == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_47 <= _pht_0_T_11;
        end else begin
          pht_0_47 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_48 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h30 == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_48 <= _pht_0_T_11;
        end else begin
          pht_0_48 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_49 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h31 == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_49 <= _pht_0_T_11;
        end else begin
          pht_0_49 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_50 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h32 == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_50 <= _pht_0_T_11;
        end else begin
          pht_0_50 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_51 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h33 == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_51 <= _pht_0_T_11;
        end else begin
          pht_0_51 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_52 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h34 == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_52 <= _pht_0_T_11;
        end else begin
          pht_0_52 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_53 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h35 == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_53 <= _pht_0_T_11;
        end else begin
          pht_0_53 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_54 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h36 == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_54 <= _pht_0_T_11;
        end else begin
          pht_0_54 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_55 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h37 == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_55 <= _pht_0_T_11;
        end else begin
          pht_0_55 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_56 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h38 == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_56 <= _pht_0_T_11;
        end else begin
          pht_0_56 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_57 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h39 == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_57 <= _pht_0_T_11;
        end else begin
          pht_0_57 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_58 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h3a == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_58 <= _pht_0_T_11;
        end else begin
          pht_0_58 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_59 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h3b == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_59 <= _pht_0_T_11;
        end else begin
          pht_0_59 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_60 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h3c == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_60 <= _pht_0_T_11;
        end else begin
          pht_0_60 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_61 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h3d == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_61 <= _pht_0_T_11;
        end else begin
          pht_0_61 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_62 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h3e == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_62 <= _pht_0_T_11;
        end else begin
          pht_0_62 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_63 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h3f == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_63 <= _pht_0_T_11;
        end else begin
          pht_0_63 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_64 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h40 == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_64 <= _pht_0_T_11;
        end else begin
          pht_0_64 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_65 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h41 == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_65 <= _pht_0_T_11;
        end else begin
          pht_0_65 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_66 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h42 == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_66 <= _pht_0_T_11;
        end else begin
          pht_0_66 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_67 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h43 == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_67 <= _pht_0_T_11;
        end else begin
          pht_0_67 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_68 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h44 == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_68 <= _pht_0_T_11;
        end else begin
          pht_0_68 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_69 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h45 == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_69 <= _pht_0_T_11;
        end else begin
          pht_0_69 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_70 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h46 == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_70 <= _pht_0_T_11;
        end else begin
          pht_0_70 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_71 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h47 == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_71 <= _pht_0_T_11;
        end else begin
          pht_0_71 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_72 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h48 == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_72 <= _pht_0_T_11;
        end else begin
          pht_0_72 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_73 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h49 == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_73 <= _pht_0_T_11;
        end else begin
          pht_0_73 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_74 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h4a == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_74 <= _pht_0_T_11;
        end else begin
          pht_0_74 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_75 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h4b == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_75 <= _pht_0_T_11;
        end else begin
          pht_0_75 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_76 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h4c == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_76 <= _pht_0_T_11;
        end else begin
          pht_0_76 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_77 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h4d == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_77 <= _pht_0_T_11;
        end else begin
          pht_0_77 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_78 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h4e == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_78 <= _pht_0_T_11;
        end else begin
          pht_0_78 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_79 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h4f == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_79 <= _pht_0_T_11;
        end else begin
          pht_0_79 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_80 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h50 == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_80 <= _pht_0_T_11;
        end else begin
          pht_0_80 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_81 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h51 == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_81 <= _pht_0_T_11;
        end else begin
          pht_0_81 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_82 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h52 == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_82 <= _pht_0_T_11;
        end else begin
          pht_0_82 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_83 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h53 == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_83 <= _pht_0_T_11;
        end else begin
          pht_0_83 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_84 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h54 == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_84 <= _pht_0_T_11;
        end else begin
          pht_0_84 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_85 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h55 == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_85 <= _pht_0_T_11;
        end else begin
          pht_0_85 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_86 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h56 == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_86 <= _pht_0_T_11;
        end else begin
          pht_0_86 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_87 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h57 == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_87 <= _pht_0_T_11;
        end else begin
          pht_0_87 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_88 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h58 == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_88 <= _pht_0_T_11;
        end else begin
          pht_0_88 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_89 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h59 == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_89 <= _pht_0_T_11;
        end else begin
          pht_0_89 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_90 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h5a == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_90 <= _pht_0_T_11;
        end else begin
          pht_0_90 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_91 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h5b == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_91 <= _pht_0_T_11;
        end else begin
          pht_0_91 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_92 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h5c == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_92 <= _pht_0_T_11;
        end else begin
          pht_0_92 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_93 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h5d == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_93 <= _pht_0_T_11;
        end else begin
          pht_0_93 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_94 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h5e == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_94 <= _pht_0_T_11;
        end else begin
          pht_0_94 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_95 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h5f == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_95 <= _pht_0_T_11;
        end else begin
          pht_0_95 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_96 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h60 == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_96 <= _pht_0_T_11;
        end else begin
          pht_0_96 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_97 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h61 == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_97 <= _pht_0_T_11;
        end else begin
          pht_0_97 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_98 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h62 == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_98 <= _pht_0_T_11;
        end else begin
          pht_0_98 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_99 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h63 == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_99 <= _pht_0_T_11;
        end else begin
          pht_0_99 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_100 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h64 == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_100 <= _pht_0_T_11;
        end else begin
          pht_0_100 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_101 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h65 == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_101 <= _pht_0_T_11;
        end else begin
          pht_0_101 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_102 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h66 == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_102 <= _pht_0_T_11;
        end else begin
          pht_0_102 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_103 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h67 == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_103 <= _pht_0_T_11;
        end else begin
          pht_0_103 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_104 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h68 == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_104 <= _pht_0_T_11;
        end else begin
          pht_0_104 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_105 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h69 == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_105 <= _pht_0_T_11;
        end else begin
          pht_0_105 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_106 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h6a == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_106 <= _pht_0_T_11;
        end else begin
          pht_0_106 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_107 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h6b == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_107 <= _pht_0_T_11;
        end else begin
          pht_0_107 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_108 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h6c == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_108 <= _pht_0_T_11;
        end else begin
          pht_0_108 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_109 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h6d == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_109 <= _pht_0_T_11;
        end else begin
          pht_0_109 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_110 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h6e == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_110 <= _pht_0_T_11;
        end else begin
          pht_0_110 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_111 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h6f == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_111 <= _pht_0_T_11;
        end else begin
          pht_0_111 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_112 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h70 == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_112 <= _pht_0_T_11;
        end else begin
          pht_0_112 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_113 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h71 == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_113 <= _pht_0_T_11;
        end else begin
          pht_0_113 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_114 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h72 == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_114 <= _pht_0_T_11;
        end else begin
          pht_0_114 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_115 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h73 == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_115 <= _pht_0_T_11;
        end else begin
          pht_0_115 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_116 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h74 == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_116 <= _pht_0_T_11;
        end else begin
          pht_0_116 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_117 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h75 == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_117 <= _pht_0_T_11;
        end else begin
          pht_0_117 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_118 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h76 == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_118 <= _pht_0_T_11;
        end else begin
          pht_0_118 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_119 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h77 == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_119 <= _pht_0_T_11;
        end else begin
          pht_0_119 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_120 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h78 == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_120 <= _pht_0_T_11;
        end else begin
          pht_0_120 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_121 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h79 == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_121 <= _pht_0_T_11;
        end else begin
          pht_0_121 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_122 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h7a == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_122 <= _pht_0_T_11;
        end else begin
          pht_0_122 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_123 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h7b == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_123 <= _pht_0_T_11;
        end else begin
          pht_0_123 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_124 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h7c == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_124 <= _pht_0_T_11;
        end else begin
          pht_0_124 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_125 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h7d == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_125 <= _pht_0_T_11;
        end else begin
          pht_0_125 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_126 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h7e == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_126 <= _pht_0_T_11;
        end else begin
          pht_0_126 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_0_127 <= 2'h1; // @[bht.scala 109:22]
    end else if (io_fire & io_takenValid) begin // @[bht.scala 161:35]
      if (7'h7f == pht1WAddr) begin // @[bht.scala 162:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_0_127 <= _pht_0_T_11;
        end else begin
          pht_0_127 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_0 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h0 == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_0 <= _pht_1_T_3;
        end else begin
          pht_1_0 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_1 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h1 == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_1 <= _pht_1_T_3;
        end else begin
          pht_1_1 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_2 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h2 == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_2 <= _pht_1_T_3;
        end else begin
          pht_1_2 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_3 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h3 == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_3 <= _pht_1_T_3;
        end else begin
          pht_1_3 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_4 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h4 == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_4 <= _pht_1_T_3;
        end else begin
          pht_1_4 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_5 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h5 == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_5 <= _pht_1_T_3;
        end else begin
          pht_1_5 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_6 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h6 == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_6 <= _pht_1_T_3;
        end else begin
          pht_1_6 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_7 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h7 == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_7 <= _pht_1_T_3;
        end else begin
          pht_1_7 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_8 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h8 == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_8 <= _pht_1_T_3;
        end else begin
          pht_1_8 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_9 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h9 == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_9 <= _pht_1_T_3;
        end else begin
          pht_1_9 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_10 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'ha == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_10 <= _pht_1_T_3;
        end else begin
          pht_1_10 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_11 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'hb == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_11 <= _pht_1_T_3;
        end else begin
          pht_1_11 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_12 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'hc == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_12 <= _pht_1_T_3;
        end else begin
          pht_1_12 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_13 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'hd == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_13 <= _pht_1_T_3;
        end else begin
          pht_1_13 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_14 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'he == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_14 <= _pht_1_T_3;
        end else begin
          pht_1_14 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_15 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'hf == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_15 <= _pht_1_T_3;
        end else begin
          pht_1_15 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_16 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h10 == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_16 <= _pht_1_T_3;
        end else begin
          pht_1_16 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_17 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h11 == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_17 <= _pht_1_T_3;
        end else begin
          pht_1_17 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_18 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h12 == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_18 <= _pht_1_T_3;
        end else begin
          pht_1_18 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_19 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h13 == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_19 <= _pht_1_T_3;
        end else begin
          pht_1_19 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_20 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h14 == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_20 <= _pht_1_T_3;
        end else begin
          pht_1_20 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_21 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h15 == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_21 <= _pht_1_T_3;
        end else begin
          pht_1_21 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_22 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h16 == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_22 <= _pht_1_T_3;
        end else begin
          pht_1_22 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_23 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h17 == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_23 <= _pht_1_T_3;
        end else begin
          pht_1_23 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_24 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h18 == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_24 <= _pht_1_T_3;
        end else begin
          pht_1_24 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_25 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h19 == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_25 <= _pht_1_T_3;
        end else begin
          pht_1_25 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_26 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h1a == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_26 <= _pht_1_T_3;
        end else begin
          pht_1_26 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_27 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h1b == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_27 <= _pht_1_T_3;
        end else begin
          pht_1_27 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_28 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h1c == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_28 <= _pht_1_T_3;
        end else begin
          pht_1_28 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_29 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h1d == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_29 <= _pht_1_T_3;
        end else begin
          pht_1_29 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_30 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h1e == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_30 <= _pht_1_T_3;
        end else begin
          pht_1_30 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_31 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h1f == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_31 <= _pht_1_T_3;
        end else begin
          pht_1_31 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_32 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h20 == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_32 <= _pht_1_T_3;
        end else begin
          pht_1_32 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_33 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h21 == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_33 <= _pht_1_T_3;
        end else begin
          pht_1_33 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_34 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h22 == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_34 <= _pht_1_T_3;
        end else begin
          pht_1_34 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_35 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h23 == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_35 <= _pht_1_T_3;
        end else begin
          pht_1_35 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_36 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h24 == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_36 <= _pht_1_T_3;
        end else begin
          pht_1_36 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_37 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h25 == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_37 <= _pht_1_T_3;
        end else begin
          pht_1_37 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_38 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h26 == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_38 <= _pht_1_T_3;
        end else begin
          pht_1_38 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_39 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h27 == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_39 <= _pht_1_T_3;
        end else begin
          pht_1_39 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_40 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h28 == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_40 <= _pht_1_T_3;
        end else begin
          pht_1_40 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_41 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h29 == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_41 <= _pht_1_T_3;
        end else begin
          pht_1_41 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_42 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h2a == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_42 <= _pht_1_T_3;
        end else begin
          pht_1_42 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_43 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h2b == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_43 <= _pht_1_T_3;
        end else begin
          pht_1_43 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_44 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h2c == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_44 <= _pht_1_T_3;
        end else begin
          pht_1_44 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_45 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h2d == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_45 <= _pht_1_T_3;
        end else begin
          pht_1_45 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_46 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h2e == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_46 <= _pht_1_T_3;
        end else begin
          pht_1_46 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_47 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h2f == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_47 <= _pht_1_T_3;
        end else begin
          pht_1_47 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_48 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h30 == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_48 <= _pht_1_T_3;
        end else begin
          pht_1_48 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_49 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h31 == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_49 <= _pht_1_T_3;
        end else begin
          pht_1_49 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_50 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h32 == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_50 <= _pht_1_T_3;
        end else begin
          pht_1_50 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_51 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h33 == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_51 <= _pht_1_T_3;
        end else begin
          pht_1_51 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_52 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h34 == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_52 <= _pht_1_T_3;
        end else begin
          pht_1_52 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_53 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h35 == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_53 <= _pht_1_T_3;
        end else begin
          pht_1_53 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_54 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h36 == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_54 <= _pht_1_T_3;
        end else begin
          pht_1_54 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_55 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h37 == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_55 <= _pht_1_T_3;
        end else begin
          pht_1_55 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_56 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h38 == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_56 <= _pht_1_T_3;
        end else begin
          pht_1_56 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_57 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h39 == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_57 <= _pht_1_T_3;
        end else begin
          pht_1_57 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_58 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h3a == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_58 <= _pht_1_T_3;
        end else begin
          pht_1_58 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_59 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h3b == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_59 <= _pht_1_T_3;
        end else begin
          pht_1_59 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_60 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h3c == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_60 <= _pht_1_T_3;
        end else begin
          pht_1_60 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_61 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h3d == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_61 <= _pht_1_T_3;
        end else begin
          pht_1_61 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_62 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h3e == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_62 <= _pht_1_T_3;
        end else begin
          pht_1_62 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_63 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h3f == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_63 <= _pht_1_T_3;
        end else begin
          pht_1_63 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_64 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h40 == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_64 <= _pht_1_T_3;
        end else begin
          pht_1_64 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_65 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h41 == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_65 <= _pht_1_T_3;
        end else begin
          pht_1_65 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_66 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h42 == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_66 <= _pht_1_T_3;
        end else begin
          pht_1_66 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_67 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h43 == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_67 <= _pht_1_T_3;
        end else begin
          pht_1_67 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_68 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h44 == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_68 <= _pht_1_T_3;
        end else begin
          pht_1_68 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_69 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h45 == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_69 <= _pht_1_T_3;
        end else begin
          pht_1_69 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_70 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h46 == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_70 <= _pht_1_T_3;
        end else begin
          pht_1_70 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_71 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h47 == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_71 <= _pht_1_T_3;
        end else begin
          pht_1_71 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_72 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h48 == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_72 <= _pht_1_T_3;
        end else begin
          pht_1_72 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_73 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h49 == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_73 <= _pht_1_T_3;
        end else begin
          pht_1_73 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_74 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h4a == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_74 <= _pht_1_T_3;
        end else begin
          pht_1_74 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_75 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h4b == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_75 <= _pht_1_T_3;
        end else begin
          pht_1_75 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_76 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h4c == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_76 <= _pht_1_T_3;
        end else begin
          pht_1_76 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_77 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h4d == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_77 <= _pht_1_T_3;
        end else begin
          pht_1_77 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_78 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h4e == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_78 <= _pht_1_T_3;
        end else begin
          pht_1_78 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_79 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h4f == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_79 <= _pht_1_T_3;
        end else begin
          pht_1_79 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_80 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h50 == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_80 <= _pht_1_T_3;
        end else begin
          pht_1_80 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_81 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h51 == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_81 <= _pht_1_T_3;
        end else begin
          pht_1_81 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_82 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h52 == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_82 <= _pht_1_T_3;
        end else begin
          pht_1_82 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_83 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h53 == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_83 <= _pht_1_T_3;
        end else begin
          pht_1_83 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_84 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h54 == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_84 <= _pht_1_T_3;
        end else begin
          pht_1_84 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_85 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h55 == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_85 <= _pht_1_T_3;
        end else begin
          pht_1_85 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_86 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h56 == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_86 <= _pht_1_T_3;
        end else begin
          pht_1_86 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_87 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h57 == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_87 <= _pht_1_T_3;
        end else begin
          pht_1_87 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_88 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h58 == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_88 <= _pht_1_T_3;
        end else begin
          pht_1_88 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_89 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h59 == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_89 <= _pht_1_T_3;
        end else begin
          pht_1_89 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_90 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h5a == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_90 <= _pht_1_T_3;
        end else begin
          pht_1_90 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_91 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h5b == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_91 <= _pht_1_T_3;
        end else begin
          pht_1_91 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_92 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h5c == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_92 <= _pht_1_T_3;
        end else begin
          pht_1_92 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_93 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h5d == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_93 <= _pht_1_T_3;
        end else begin
          pht_1_93 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_94 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h5e == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_94 <= _pht_1_T_3;
        end else begin
          pht_1_94 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_95 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h5f == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_95 <= _pht_1_T_3;
        end else begin
          pht_1_95 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_96 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h60 == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_96 <= _pht_1_T_3;
        end else begin
          pht_1_96 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_97 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h61 == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_97 <= _pht_1_T_3;
        end else begin
          pht_1_97 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_98 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h62 == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_98 <= _pht_1_T_3;
        end else begin
          pht_1_98 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_99 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h63 == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_99 <= _pht_1_T_3;
        end else begin
          pht_1_99 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_100 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h64 == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_100 <= _pht_1_T_3;
        end else begin
          pht_1_100 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_101 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h65 == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_101 <= _pht_1_T_3;
        end else begin
          pht_1_101 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_102 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h66 == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_102 <= _pht_1_T_3;
        end else begin
          pht_1_102 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_103 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h67 == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_103 <= _pht_1_T_3;
        end else begin
          pht_1_103 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_104 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h68 == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_104 <= _pht_1_T_3;
        end else begin
          pht_1_104 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_105 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h69 == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_105 <= _pht_1_T_3;
        end else begin
          pht_1_105 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_106 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h6a == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_106 <= _pht_1_T_3;
        end else begin
          pht_1_106 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_107 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h6b == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_107 <= _pht_1_T_3;
        end else begin
          pht_1_107 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_108 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h6c == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_108 <= _pht_1_T_3;
        end else begin
          pht_1_108 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_109 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h6d == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_109 <= _pht_1_T_3;
        end else begin
          pht_1_109 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_110 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h6e == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_110 <= _pht_1_T_3;
        end else begin
          pht_1_110 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_111 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h6f == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_111 <= _pht_1_T_3;
        end else begin
          pht_1_111 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_112 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h70 == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_112 <= _pht_1_T_3;
        end else begin
          pht_1_112 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_113 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h71 == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_113 <= _pht_1_T_3;
        end else begin
          pht_1_113 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_114 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h72 == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_114 <= _pht_1_T_3;
        end else begin
          pht_1_114 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_115 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h73 == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_115 <= _pht_1_T_3;
        end else begin
          pht_1_115 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_116 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h74 == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_116 <= _pht_1_T_3;
        end else begin
          pht_1_116 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_117 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h75 == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_117 <= _pht_1_T_3;
        end else begin
          pht_1_117 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_118 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h76 == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_118 <= _pht_1_T_3;
        end else begin
          pht_1_118 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_119 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h77 == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_119 <= _pht_1_T_3;
        end else begin
          pht_1_119 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_120 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h78 == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_120 <= _pht_1_T_3;
        end else begin
          pht_1_120 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_121 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h79 == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_121 <= _pht_1_T_3;
        end else begin
          pht_1_121 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_122 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h7a == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_122 <= _pht_1_T_3;
        end else begin
          pht_1_122 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_123 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h7b == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_123 <= _pht_1_T_3;
        end else begin
          pht_1_123 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_124 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h7c == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_124 <= _pht_1_T_3;
        end else begin
          pht_1_124 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_125 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h7d == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_125 <= _pht_1_T_3;
        end else begin
          pht_1_125 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_126 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h7e == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_126 <= _pht_1_T_3;
        end else begin
          pht_1_126 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_1_127 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 171:35]
      if (7'h7f == pht1WAddr) begin // @[bht.scala 172:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_127 <= _pht_1_T_3;
        end else begin
          pht_1_127 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_0 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h0 == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_0 <= _pht_1_T_3;
        end else begin
          pht_2_0 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_1 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h1 == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_1 <= _pht_1_T_3;
        end else begin
          pht_2_1 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_2 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h2 == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_2 <= _pht_1_T_3;
        end else begin
          pht_2_2 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_3 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h3 == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_3 <= _pht_1_T_3;
        end else begin
          pht_2_3 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_4 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h4 == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_4 <= _pht_1_T_3;
        end else begin
          pht_2_4 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_5 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h5 == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_5 <= _pht_1_T_3;
        end else begin
          pht_2_5 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_6 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h6 == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_6 <= _pht_1_T_3;
        end else begin
          pht_2_6 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_7 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h7 == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_7 <= _pht_1_T_3;
        end else begin
          pht_2_7 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_8 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h8 == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_8 <= _pht_1_T_3;
        end else begin
          pht_2_8 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_9 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h9 == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_9 <= _pht_1_T_3;
        end else begin
          pht_2_9 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_10 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'ha == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_10 <= _pht_1_T_3;
        end else begin
          pht_2_10 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_11 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'hb == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_11 <= _pht_1_T_3;
        end else begin
          pht_2_11 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_12 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'hc == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_12 <= _pht_1_T_3;
        end else begin
          pht_2_12 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_13 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'hd == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_13 <= _pht_1_T_3;
        end else begin
          pht_2_13 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_14 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'he == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_14 <= _pht_1_T_3;
        end else begin
          pht_2_14 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_15 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'hf == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_15 <= _pht_1_T_3;
        end else begin
          pht_2_15 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_16 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h10 == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_16 <= _pht_1_T_3;
        end else begin
          pht_2_16 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_17 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h11 == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_17 <= _pht_1_T_3;
        end else begin
          pht_2_17 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_18 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h12 == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_18 <= _pht_1_T_3;
        end else begin
          pht_2_18 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_19 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h13 == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_19 <= _pht_1_T_3;
        end else begin
          pht_2_19 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_20 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h14 == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_20 <= _pht_1_T_3;
        end else begin
          pht_2_20 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_21 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h15 == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_21 <= _pht_1_T_3;
        end else begin
          pht_2_21 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_22 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h16 == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_22 <= _pht_1_T_3;
        end else begin
          pht_2_22 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_23 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h17 == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_23 <= _pht_1_T_3;
        end else begin
          pht_2_23 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_24 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h18 == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_24 <= _pht_1_T_3;
        end else begin
          pht_2_24 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_25 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h19 == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_25 <= _pht_1_T_3;
        end else begin
          pht_2_25 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_26 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h1a == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_26 <= _pht_1_T_3;
        end else begin
          pht_2_26 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_27 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h1b == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_27 <= _pht_1_T_3;
        end else begin
          pht_2_27 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_28 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h1c == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_28 <= _pht_1_T_3;
        end else begin
          pht_2_28 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_29 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h1d == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_29 <= _pht_1_T_3;
        end else begin
          pht_2_29 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_30 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h1e == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_30 <= _pht_1_T_3;
        end else begin
          pht_2_30 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_31 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h1f == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_31 <= _pht_1_T_3;
        end else begin
          pht_2_31 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_32 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h20 == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_32 <= _pht_1_T_3;
        end else begin
          pht_2_32 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_33 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h21 == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_33 <= _pht_1_T_3;
        end else begin
          pht_2_33 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_34 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h22 == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_34 <= _pht_1_T_3;
        end else begin
          pht_2_34 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_35 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h23 == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_35 <= _pht_1_T_3;
        end else begin
          pht_2_35 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_36 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h24 == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_36 <= _pht_1_T_3;
        end else begin
          pht_2_36 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_37 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h25 == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_37 <= _pht_1_T_3;
        end else begin
          pht_2_37 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_38 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h26 == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_38 <= _pht_1_T_3;
        end else begin
          pht_2_38 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_39 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h27 == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_39 <= _pht_1_T_3;
        end else begin
          pht_2_39 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_40 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h28 == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_40 <= _pht_1_T_3;
        end else begin
          pht_2_40 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_41 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h29 == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_41 <= _pht_1_T_3;
        end else begin
          pht_2_41 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_42 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h2a == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_42 <= _pht_1_T_3;
        end else begin
          pht_2_42 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_43 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h2b == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_43 <= _pht_1_T_3;
        end else begin
          pht_2_43 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_44 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h2c == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_44 <= _pht_1_T_3;
        end else begin
          pht_2_44 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_45 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h2d == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_45 <= _pht_1_T_3;
        end else begin
          pht_2_45 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_46 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h2e == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_46 <= _pht_1_T_3;
        end else begin
          pht_2_46 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_47 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h2f == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_47 <= _pht_1_T_3;
        end else begin
          pht_2_47 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_48 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h30 == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_48 <= _pht_1_T_3;
        end else begin
          pht_2_48 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_49 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h31 == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_49 <= _pht_1_T_3;
        end else begin
          pht_2_49 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_50 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h32 == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_50 <= _pht_1_T_3;
        end else begin
          pht_2_50 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_51 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h33 == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_51 <= _pht_1_T_3;
        end else begin
          pht_2_51 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_52 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h34 == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_52 <= _pht_1_T_3;
        end else begin
          pht_2_52 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_53 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h35 == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_53 <= _pht_1_T_3;
        end else begin
          pht_2_53 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_54 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h36 == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_54 <= _pht_1_T_3;
        end else begin
          pht_2_54 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_55 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h37 == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_55 <= _pht_1_T_3;
        end else begin
          pht_2_55 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_56 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h38 == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_56 <= _pht_1_T_3;
        end else begin
          pht_2_56 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_57 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h39 == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_57 <= _pht_1_T_3;
        end else begin
          pht_2_57 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_58 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h3a == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_58 <= _pht_1_T_3;
        end else begin
          pht_2_58 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_59 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h3b == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_59 <= _pht_1_T_3;
        end else begin
          pht_2_59 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_60 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h3c == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_60 <= _pht_1_T_3;
        end else begin
          pht_2_60 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_61 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h3d == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_61 <= _pht_1_T_3;
        end else begin
          pht_2_61 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_62 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h3e == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_62 <= _pht_1_T_3;
        end else begin
          pht_2_62 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_63 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h3f == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_63 <= _pht_1_T_3;
        end else begin
          pht_2_63 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_64 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h40 == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_64 <= _pht_1_T_3;
        end else begin
          pht_2_64 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_65 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h41 == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_65 <= _pht_1_T_3;
        end else begin
          pht_2_65 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_66 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h42 == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_66 <= _pht_1_T_3;
        end else begin
          pht_2_66 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_67 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h43 == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_67 <= _pht_1_T_3;
        end else begin
          pht_2_67 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_68 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h44 == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_68 <= _pht_1_T_3;
        end else begin
          pht_2_68 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_69 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h45 == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_69 <= _pht_1_T_3;
        end else begin
          pht_2_69 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_70 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h46 == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_70 <= _pht_1_T_3;
        end else begin
          pht_2_70 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_71 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h47 == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_71 <= _pht_1_T_3;
        end else begin
          pht_2_71 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_72 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h48 == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_72 <= _pht_1_T_3;
        end else begin
          pht_2_72 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_73 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h49 == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_73 <= _pht_1_T_3;
        end else begin
          pht_2_73 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_74 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h4a == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_74 <= _pht_1_T_3;
        end else begin
          pht_2_74 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_75 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h4b == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_75 <= _pht_1_T_3;
        end else begin
          pht_2_75 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_76 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h4c == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_76 <= _pht_1_T_3;
        end else begin
          pht_2_76 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_77 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h4d == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_77 <= _pht_1_T_3;
        end else begin
          pht_2_77 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_78 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h4e == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_78 <= _pht_1_T_3;
        end else begin
          pht_2_78 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_79 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h4f == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_79 <= _pht_1_T_3;
        end else begin
          pht_2_79 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_80 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h50 == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_80 <= _pht_1_T_3;
        end else begin
          pht_2_80 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_81 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h51 == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_81 <= _pht_1_T_3;
        end else begin
          pht_2_81 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_82 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h52 == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_82 <= _pht_1_T_3;
        end else begin
          pht_2_82 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_83 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h53 == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_83 <= _pht_1_T_3;
        end else begin
          pht_2_83 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_84 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h54 == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_84 <= _pht_1_T_3;
        end else begin
          pht_2_84 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_85 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h55 == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_85 <= _pht_1_T_3;
        end else begin
          pht_2_85 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_86 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h56 == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_86 <= _pht_1_T_3;
        end else begin
          pht_2_86 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_87 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h57 == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_87 <= _pht_1_T_3;
        end else begin
          pht_2_87 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_88 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h58 == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_88 <= _pht_1_T_3;
        end else begin
          pht_2_88 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_89 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h59 == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_89 <= _pht_1_T_3;
        end else begin
          pht_2_89 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_90 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h5a == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_90 <= _pht_1_T_3;
        end else begin
          pht_2_90 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_91 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h5b == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_91 <= _pht_1_T_3;
        end else begin
          pht_2_91 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_92 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h5c == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_92 <= _pht_1_T_3;
        end else begin
          pht_2_92 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_93 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h5d == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_93 <= _pht_1_T_3;
        end else begin
          pht_2_93 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_94 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h5e == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_94 <= _pht_1_T_3;
        end else begin
          pht_2_94 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_95 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h5f == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_95 <= _pht_1_T_3;
        end else begin
          pht_2_95 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_96 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h60 == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_96 <= _pht_1_T_3;
        end else begin
          pht_2_96 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_97 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h61 == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_97 <= _pht_1_T_3;
        end else begin
          pht_2_97 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_98 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h62 == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_98 <= _pht_1_T_3;
        end else begin
          pht_2_98 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_99 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h63 == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_99 <= _pht_1_T_3;
        end else begin
          pht_2_99 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_100 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h64 == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_100 <= _pht_1_T_3;
        end else begin
          pht_2_100 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_101 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h65 == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_101 <= _pht_1_T_3;
        end else begin
          pht_2_101 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_102 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h66 == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_102 <= _pht_1_T_3;
        end else begin
          pht_2_102 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_103 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h67 == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_103 <= _pht_1_T_3;
        end else begin
          pht_2_103 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_104 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h68 == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_104 <= _pht_1_T_3;
        end else begin
          pht_2_104 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_105 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h69 == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_105 <= _pht_1_T_3;
        end else begin
          pht_2_105 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_106 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h6a == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_106 <= _pht_1_T_3;
        end else begin
          pht_2_106 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_107 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h6b == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_107 <= _pht_1_T_3;
        end else begin
          pht_2_107 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_108 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h6c == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_108 <= _pht_1_T_3;
        end else begin
          pht_2_108 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_109 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h6d == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_109 <= _pht_1_T_3;
        end else begin
          pht_2_109 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_110 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h6e == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_110 <= _pht_1_T_3;
        end else begin
          pht_2_110 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_111 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h6f == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_111 <= _pht_1_T_3;
        end else begin
          pht_2_111 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_112 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h70 == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_112 <= _pht_1_T_3;
        end else begin
          pht_2_112 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_113 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h71 == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_113 <= _pht_1_T_3;
        end else begin
          pht_2_113 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_114 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h72 == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_114 <= _pht_1_T_3;
        end else begin
          pht_2_114 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_115 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h73 == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_115 <= _pht_1_T_3;
        end else begin
          pht_2_115 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_116 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h74 == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_116 <= _pht_1_T_3;
        end else begin
          pht_2_116 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_117 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h75 == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_117 <= _pht_1_T_3;
        end else begin
          pht_2_117 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_118 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h76 == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_118 <= _pht_1_T_3;
        end else begin
          pht_2_118 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_119 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h77 == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_119 <= _pht_1_T_3;
        end else begin
          pht_2_119 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_120 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h78 == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_120 <= _pht_1_T_3;
        end else begin
          pht_2_120 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_121 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h79 == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_121 <= _pht_1_T_3;
        end else begin
          pht_2_121 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_122 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h7a == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_122 <= _pht_1_T_3;
        end else begin
          pht_2_122 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_123 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h7b == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_123 <= _pht_1_T_3;
        end else begin
          pht_2_123 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_124 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h7c == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_124 <= _pht_1_T_3;
        end else begin
          pht_2_124 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_125 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h7d == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_125 <= _pht_1_T_3;
        end else begin
          pht_2_125 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_126 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h7e == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_126 <= _pht_1_T_3;
        end else begin
          pht_2_126 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 109:22]
      pht_2_127 <= 2'h1; // @[bht.scala 109:22]
    end else if (_T) begin // @[bht.scala 179:35]
      if (7'h7f == pht2WAddr) begin // @[bht.scala 180:25]
        if (2'h3 == _GEN_1279) begin // @[Mux.scala 81:58]
          pht_2_127 <= _pht_1_T_3;
        end else begin
          pht_2_127 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_0 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_0 <= _GEN_2433;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_1 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_1 <= _GEN_2434;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_2 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_2 <= _GEN_2435;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_3 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_3 <= _GEN_2436;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_4 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_4 <= _GEN_2437;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_5 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_5 <= _GEN_2438;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_6 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_6 <= _GEN_2439;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_7 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_7 <= _GEN_2440;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_8 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_8 <= _GEN_2441;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_9 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_9 <= _GEN_2442;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_10 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_10 <= _GEN_2443;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_11 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_11 <= _GEN_2444;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_12 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_12 <= _GEN_2445;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_13 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_13 <= _GEN_2446;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_14 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_14 <= _GEN_2447;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_15 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_15 <= _GEN_2448;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_16 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_16 <= _GEN_2449;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_17 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_17 <= _GEN_2450;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_18 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_18 <= _GEN_2451;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_19 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_19 <= _GEN_2452;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_20 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_20 <= _GEN_2453;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_21 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_21 <= _GEN_2454;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_22 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_22 <= _GEN_2455;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_23 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_23 <= _GEN_2456;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_24 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_24 <= _GEN_2457;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_25 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_25 <= _GEN_2458;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_26 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_26 <= _GEN_2459;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_27 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_27 <= _GEN_2460;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_28 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_28 <= _GEN_2461;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_29 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_29 <= _GEN_2462;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_30 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_30 <= _GEN_2463;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_31 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_31 <= _GEN_2464;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_32 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_32 <= _GEN_2465;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_33 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_33 <= _GEN_2466;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_34 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_34 <= _GEN_2467;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_35 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_35 <= _GEN_2468;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_36 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_36 <= _GEN_2469;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_37 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_37 <= _GEN_2470;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_38 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_38 <= _GEN_2471;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_39 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_39 <= _GEN_2472;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_40 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_40 <= _GEN_2473;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_41 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_41 <= _GEN_2474;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_42 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_42 <= _GEN_2475;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_43 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_43 <= _GEN_2476;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_44 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_44 <= _GEN_2477;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_45 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_45 <= _GEN_2478;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_46 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_46 <= _GEN_2479;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_47 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_47 <= _GEN_2480;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_48 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_48 <= _GEN_2481;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_49 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_49 <= _GEN_2482;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_50 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_50 <= _GEN_2483;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_51 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_51 <= _GEN_2484;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_52 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_52 <= _GEN_2485;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_53 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_53 <= _GEN_2486;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_54 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_54 <= _GEN_2487;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_55 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_55 <= _GEN_2488;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_56 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_56 <= _GEN_2489;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_57 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_57 <= _GEN_2490;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_58 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_58 <= _GEN_2491;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_59 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_59 <= _GEN_2492;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_60 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_60 <= _GEN_2493;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_61 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_61 <= _GEN_2494;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_62 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_62 <= _GEN_2495;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_63 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_63 <= _GEN_2496;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_64 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_64 <= _GEN_2497;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_65 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_65 <= _GEN_2498;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_66 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_66 <= _GEN_2499;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_67 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_67 <= _GEN_2500;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_68 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_68 <= _GEN_2501;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_69 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_69 <= _GEN_2502;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_70 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_70 <= _GEN_2503;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_71 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_71 <= _GEN_2504;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_72 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_72 <= _GEN_2505;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_73 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_73 <= _GEN_2506;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_74 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_74 <= _GEN_2507;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_75 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_75 <= _GEN_2508;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_76 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_76 <= _GEN_2509;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_77 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_77 <= _GEN_2510;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_78 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_78 <= _GEN_2511;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_79 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_79 <= _GEN_2512;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_80 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_80 <= _GEN_2513;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_81 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_81 <= _GEN_2514;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_82 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_82 <= _GEN_2515;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_83 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_83 <= _GEN_2516;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_84 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_84 <= _GEN_2517;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_85 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_85 <= _GEN_2518;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_86 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_86 <= _GEN_2519;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_87 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_87 <= _GEN_2520;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_88 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_88 <= _GEN_2521;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_89 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_89 <= _GEN_2522;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_90 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_90 <= _GEN_2523;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_91 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_91 <= _GEN_2524;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_92 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_92 <= _GEN_2525;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_93 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_93 <= _GEN_2526;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_94 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_94 <= _GEN_2527;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_95 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_95 <= _GEN_2528;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_96 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_96 <= _GEN_2529;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_97 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_97 <= _GEN_2530;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_98 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_98 <= _GEN_2531;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_99 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_99 <= _GEN_2532;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_100 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_100 <= _GEN_2533;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_101 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_101 <= _GEN_2534;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_102 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_102 <= _GEN_2535;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_103 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_103 <= _GEN_2536;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_104 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_104 <= _GEN_2537;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_105 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_105 <= _GEN_2538;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_106 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_106 <= _GEN_2539;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_107 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_107 <= _GEN_2540;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_108 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_108 <= _GEN_2541;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_109 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_109 <= _GEN_2542;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_110 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_110 <= _GEN_2543;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_111 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_111 <= _GEN_2544;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_112 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_112 <= _GEN_2545;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_113 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_113 <= _GEN_2546;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_114 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_114 <= _GEN_2547;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_115 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_115 <= _GEN_2548;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_116 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_116 <= _GEN_2549;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_117 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_117 <= _GEN_2550;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_118 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_118 <= _GEN_2551;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_119 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_119 <= _GEN_2552;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_120 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_120 <= _GEN_2553;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_121 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_121 <= _GEN_2554;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_122 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_122 <= _GEN_2555;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_123 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_123 <= _GEN_2556;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_124 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_124 <= _GEN_2557;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_125 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_125 <= _GEN_2558;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_126 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_126 <= _GEN_2559;
    end
    if (reset) begin // @[bht.scala 112:23]
      btbV_127 <= 1'h0; // @[bht.scala 112:23]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      btbV_127 <= _GEN_2560;
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_0 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h0 == upIndex) begin // @[bht.scala 199:21]
        btbTag_0 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_1 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h1 == upIndex) begin // @[bht.scala 199:21]
        btbTag_1 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_2 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h2 == upIndex) begin // @[bht.scala 199:21]
        btbTag_2 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_3 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h3 == upIndex) begin // @[bht.scala 199:21]
        btbTag_3 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_4 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h4 == upIndex) begin // @[bht.scala 199:21]
        btbTag_4 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_5 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h5 == upIndex) begin // @[bht.scala 199:21]
        btbTag_5 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_6 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h6 == upIndex) begin // @[bht.scala 199:21]
        btbTag_6 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_7 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h7 == upIndex) begin // @[bht.scala 199:21]
        btbTag_7 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_8 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h8 == upIndex) begin // @[bht.scala 199:21]
        btbTag_8 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_9 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h9 == upIndex) begin // @[bht.scala 199:21]
        btbTag_9 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_10 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'ha == upIndex) begin // @[bht.scala 199:21]
        btbTag_10 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_11 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'hb == upIndex) begin // @[bht.scala 199:21]
        btbTag_11 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_12 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'hc == upIndex) begin // @[bht.scala 199:21]
        btbTag_12 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_13 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'hd == upIndex) begin // @[bht.scala 199:21]
        btbTag_13 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_14 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'he == upIndex) begin // @[bht.scala 199:21]
        btbTag_14 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_15 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'hf == upIndex) begin // @[bht.scala 199:21]
        btbTag_15 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_16 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h10 == upIndex) begin // @[bht.scala 199:21]
        btbTag_16 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_17 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h11 == upIndex) begin // @[bht.scala 199:21]
        btbTag_17 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_18 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h12 == upIndex) begin // @[bht.scala 199:21]
        btbTag_18 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_19 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h13 == upIndex) begin // @[bht.scala 199:21]
        btbTag_19 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_20 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h14 == upIndex) begin // @[bht.scala 199:21]
        btbTag_20 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_21 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h15 == upIndex) begin // @[bht.scala 199:21]
        btbTag_21 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_22 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h16 == upIndex) begin // @[bht.scala 199:21]
        btbTag_22 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_23 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h17 == upIndex) begin // @[bht.scala 199:21]
        btbTag_23 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_24 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h18 == upIndex) begin // @[bht.scala 199:21]
        btbTag_24 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_25 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h19 == upIndex) begin // @[bht.scala 199:21]
        btbTag_25 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_26 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h1a == upIndex) begin // @[bht.scala 199:21]
        btbTag_26 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_27 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h1b == upIndex) begin // @[bht.scala 199:21]
        btbTag_27 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_28 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h1c == upIndex) begin // @[bht.scala 199:21]
        btbTag_28 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_29 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h1d == upIndex) begin // @[bht.scala 199:21]
        btbTag_29 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_30 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h1e == upIndex) begin // @[bht.scala 199:21]
        btbTag_30 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_31 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h1f == upIndex) begin // @[bht.scala 199:21]
        btbTag_31 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_32 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h20 == upIndex) begin // @[bht.scala 199:21]
        btbTag_32 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_33 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h21 == upIndex) begin // @[bht.scala 199:21]
        btbTag_33 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_34 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h22 == upIndex) begin // @[bht.scala 199:21]
        btbTag_34 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_35 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h23 == upIndex) begin // @[bht.scala 199:21]
        btbTag_35 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_36 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h24 == upIndex) begin // @[bht.scala 199:21]
        btbTag_36 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_37 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h25 == upIndex) begin // @[bht.scala 199:21]
        btbTag_37 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_38 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h26 == upIndex) begin // @[bht.scala 199:21]
        btbTag_38 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_39 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h27 == upIndex) begin // @[bht.scala 199:21]
        btbTag_39 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_40 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h28 == upIndex) begin // @[bht.scala 199:21]
        btbTag_40 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_41 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h29 == upIndex) begin // @[bht.scala 199:21]
        btbTag_41 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_42 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h2a == upIndex) begin // @[bht.scala 199:21]
        btbTag_42 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_43 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h2b == upIndex) begin // @[bht.scala 199:21]
        btbTag_43 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_44 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h2c == upIndex) begin // @[bht.scala 199:21]
        btbTag_44 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_45 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h2d == upIndex) begin // @[bht.scala 199:21]
        btbTag_45 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_46 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h2e == upIndex) begin // @[bht.scala 199:21]
        btbTag_46 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_47 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h2f == upIndex) begin // @[bht.scala 199:21]
        btbTag_47 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_48 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h30 == upIndex) begin // @[bht.scala 199:21]
        btbTag_48 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_49 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h31 == upIndex) begin // @[bht.scala 199:21]
        btbTag_49 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_50 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h32 == upIndex) begin // @[bht.scala 199:21]
        btbTag_50 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_51 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h33 == upIndex) begin // @[bht.scala 199:21]
        btbTag_51 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_52 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h34 == upIndex) begin // @[bht.scala 199:21]
        btbTag_52 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_53 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h35 == upIndex) begin // @[bht.scala 199:21]
        btbTag_53 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_54 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h36 == upIndex) begin // @[bht.scala 199:21]
        btbTag_54 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_55 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h37 == upIndex) begin // @[bht.scala 199:21]
        btbTag_55 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_56 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h38 == upIndex) begin // @[bht.scala 199:21]
        btbTag_56 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_57 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h39 == upIndex) begin // @[bht.scala 199:21]
        btbTag_57 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_58 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h3a == upIndex) begin // @[bht.scala 199:21]
        btbTag_58 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_59 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h3b == upIndex) begin // @[bht.scala 199:21]
        btbTag_59 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_60 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h3c == upIndex) begin // @[bht.scala 199:21]
        btbTag_60 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_61 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h3d == upIndex) begin // @[bht.scala 199:21]
        btbTag_61 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_62 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h3e == upIndex) begin // @[bht.scala 199:21]
        btbTag_62 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_63 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h3f == upIndex) begin // @[bht.scala 199:21]
        btbTag_63 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_64 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h40 == upIndex) begin // @[bht.scala 199:21]
        btbTag_64 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_65 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h41 == upIndex) begin // @[bht.scala 199:21]
        btbTag_65 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_66 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h42 == upIndex) begin // @[bht.scala 199:21]
        btbTag_66 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_67 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h43 == upIndex) begin // @[bht.scala 199:21]
        btbTag_67 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_68 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h44 == upIndex) begin // @[bht.scala 199:21]
        btbTag_68 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_69 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h45 == upIndex) begin // @[bht.scala 199:21]
        btbTag_69 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_70 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h46 == upIndex) begin // @[bht.scala 199:21]
        btbTag_70 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_71 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h47 == upIndex) begin // @[bht.scala 199:21]
        btbTag_71 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_72 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h48 == upIndex) begin // @[bht.scala 199:21]
        btbTag_72 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_73 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h49 == upIndex) begin // @[bht.scala 199:21]
        btbTag_73 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_74 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h4a == upIndex) begin // @[bht.scala 199:21]
        btbTag_74 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_75 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h4b == upIndex) begin // @[bht.scala 199:21]
        btbTag_75 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_76 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h4c == upIndex) begin // @[bht.scala 199:21]
        btbTag_76 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_77 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h4d == upIndex) begin // @[bht.scala 199:21]
        btbTag_77 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_78 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h4e == upIndex) begin // @[bht.scala 199:21]
        btbTag_78 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_79 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h4f == upIndex) begin // @[bht.scala 199:21]
        btbTag_79 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_80 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h50 == upIndex) begin // @[bht.scala 199:21]
        btbTag_80 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_81 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h51 == upIndex) begin // @[bht.scala 199:21]
        btbTag_81 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_82 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h52 == upIndex) begin // @[bht.scala 199:21]
        btbTag_82 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_83 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h53 == upIndex) begin // @[bht.scala 199:21]
        btbTag_83 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_84 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h54 == upIndex) begin // @[bht.scala 199:21]
        btbTag_84 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_85 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h55 == upIndex) begin // @[bht.scala 199:21]
        btbTag_85 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_86 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h56 == upIndex) begin // @[bht.scala 199:21]
        btbTag_86 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_87 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h57 == upIndex) begin // @[bht.scala 199:21]
        btbTag_87 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_88 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h58 == upIndex) begin // @[bht.scala 199:21]
        btbTag_88 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_89 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h59 == upIndex) begin // @[bht.scala 199:21]
        btbTag_89 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_90 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h5a == upIndex) begin // @[bht.scala 199:21]
        btbTag_90 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_91 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h5b == upIndex) begin // @[bht.scala 199:21]
        btbTag_91 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_92 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h5c == upIndex) begin // @[bht.scala 199:21]
        btbTag_92 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_93 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h5d == upIndex) begin // @[bht.scala 199:21]
        btbTag_93 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_94 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h5e == upIndex) begin // @[bht.scala 199:21]
        btbTag_94 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_95 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h5f == upIndex) begin // @[bht.scala 199:21]
        btbTag_95 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_96 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h60 == upIndex) begin // @[bht.scala 199:21]
        btbTag_96 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_97 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h61 == upIndex) begin // @[bht.scala 199:21]
        btbTag_97 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_98 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h62 == upIndex) begin // @[bht.scala 199:21]
        btbTag_98 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_99 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h63 == upIndex) begin // @[bht.scala 199:21]
        btbTag_99 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_100 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h64 == upIndex) begin // @[bht.scala 199:21]
        btbTag_100 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_101 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h65 == upIndex) begin // @[bht.scala 199:21]
        btbTag_101 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_102 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h66 == upIndex) begin // @[bht.scala 199:21]
        btbTag_102 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_103 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h67 == upIndex) begin // @[bht.scala 199:21]
        btbTag_103 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_104 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h68 == upIndex) begin // @[bht.scala 199:21]
        btbTag_104 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_105 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h69 == upIndex) begin // @[bht.scala 199:21]
        btbTag_105 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_106 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h6a == upIndex) begin // @[bht.scala 199:21]
        btbTag_106 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_107 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h6b == upIndex) begin // @[bht.scala 199:21]
        btbTag_107 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_108 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h6c == upIndex) begin // @[bht.scala 199:21]
        btbTag_108 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_109 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h6d == upIndex) begin // @[bht.scala 199:21]
        btbTag_109 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_110 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h6e == upIndex) begin // @[bht.scala 199:21]
        btbTag_110 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_111 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h6f == upIndex) begin // @[bht.scala 199:21]
        btbTag_111 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_112 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h70 == upIndex) begin // @[bht.scala 199:21]
        btbTag_112 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_113 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h71 == upIndex) begin // @[bht.scala 199:21]
        btbTag_113 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_114 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h72 == upIndex) begin // @[bht.scala 199:21]
        btbTag_114 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_115 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h73 == upIndex) begin // @[bht.scala 199:21]
        btbTag_115 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_116 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h74 == upIndex) begin // @[bht.scala 199:21]
        btbTag_116 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_117 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h75 == upIndex) begin // @[bht.scala 199:21]
        btbTag_117 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_118 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h76 == upIndex) begin // @[bht.scala 199:21]
        btbTag_118 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_119 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h77 == upIndex) begin // @[bht.scala 199:21]
        btbTag_119 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_120 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h78 == upIndex) begin // @[bht.scala 199:21]
        btbTag_120 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_121 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h79 == upIndex) begin // @[bht.scala 199:21]
        btbTag_121 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_122 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h7a == upIndex) begin // @[bht.scala 199:21]
        btbTag_122 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_123 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h7b == upIndex) begin // @[bht.scala 199:21]
        btbTag_123 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_124 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h7c == upIndex) begin // @[bht.scala 199:21]
        btbTag_124 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_125 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h7d == upIndex) begin // @[bht.scala 199:21]
        btbTag_125 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_126 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h7e == upIndex) begin // @[bht.scala 199:21]
        btbTag_126 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 113:25]
      btbTag_127 <= 7'h0; // @[bht.scala 113:25]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h7f == upIndex) begin // @[bht.scala 199:21]
        btbTag_127 <= bhtWAddr; // @[bht.scala 199:21]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_0 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h0 == upIndex) begin // @[bht.scala 200:22]
        btbMeta_0 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_1 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h1 == upIndex) begin // @[bht.scala 200:22]
        btbMeta_1 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_2 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h2 == upIndex) begin // @[bht.scala 200:22]
        btbMeta_2 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_3 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h3 == upIndex) begin // @[bht.scala 200:22]
        btbMeta_3 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_4 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h4 == upIndex) begin // @[bht.scala 200:22]
        btbMeta_4 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_5 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h5 == upIndex) begin // @[bht.scala 200:22]
        btbMeta_5 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_6 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h6 == upIndex) begin // @[bht.scala 200:22]
        btbMeta_6 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_7 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h7 == upIndex) begin // @[bht.scala 200:22]
        btbMeta_7 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_8 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h8 == upIndex) begin // @[bht.scala 200:22]
        btbMeta_8 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_9 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h9 == upIndex) begin // @[bht.scala 200:22]
        btbMeta_9 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_10 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'ha == upIndex) begin // @[bht.scala 200:22]
        btbMeta_10 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_11 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'hb == upIndex) begin // @[bht.scala 200:22]
        btbMeta_11 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_12 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'hc == upIndex) begin // @[bht.scala 200:22]
        btbMeta_12 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_13 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'hd == upIndex) begin // @[bht.scala 200:22]
        btbMeta_13 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_14 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'he == upIndex) begin // @[bht.scala 200:22]
        btbMeta_14 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_15 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'hf == upIndex) begin // @[bht.scala 200:22]
        btbMeta_15 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_16 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h10 == upIndex) begin // @[bht.scala 200:22]
        btbMeta_16 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_17 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h11 == upIndex) begin // @[bht.scala 200:22]
        btbMeta_17 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_18 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h12 == upIndex) begin // @[bht.scala 200:22]
        btbMeta_18 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_19 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h13 == upIndex) begin // @[bht.scala 200:22]
        btbMeta_19 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_20 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h14 == upIndex) begin // @[bht.scala 200:22]
        btbMeta_20 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_21 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h15 == upIndex) begin // @[bht.scala 200:22]
        btbMeta_21 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_22 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h16 == upIndex) begin // @[bht.scala 200:22]
        btbMeta_22 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_23 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h17 == upIndex) begin // @[bht.scala 200:22]
        btbMeta_23 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_24 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h18 == upIndex) begin // @[bht.scala 200:22]
        btbMeta_24 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_25 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h19 == upIndex) begin // @[bht.scala 200:22]
        btbMeta_25 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_26 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h1a == upIndex) begin // @[bht.scala 200:22]
        btbMeta_26 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_27 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h1b == upIndex) begin // @[bht.scala 200:22]
        btbMeta_27 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_28 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h1c == upIndex) begin // @[bht.scala 200:22]
        btbMeta_28 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_29 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h1d == upIndex) begin // @[bht.scala 200:22]
        btbMeta_29 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_30 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h1e == upIndex) begin // @[bht.scala 200:22]
        btbMeta_30 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_31 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h1f == upIndex) begin // @[bht.scala 200:22]
        btbMeta_31 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_32 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h20 == upIndex) begin // @[bht.scala 200:22]
        btbMeta_32 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_33 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h21 == upIndex) begin // @[bht.scala 200:22]
        btbMeta_33 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_34 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h22 == upIndex) begin // @[bht.scala 200:22]
        btbMeta_34 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_35 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h23 == upIndex) begin // @[bht.scala 200:22]
        btbMeta_35 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_36 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h24 == upIndex) begin // @[bht.scala 200:22]
        btbMeta_36 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_37 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h25 == upIndex) begin // @[bht.scala 200:22]
        btbMeta_37 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_38 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h26 == upIndex) begin // @[bht.scala 200:22]
        btbMeta_38 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_39 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h27 == upIndex) begin // @[bht.scala 200:22]
        btbMeta_39 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_40 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h28 == upIndex) begin // @[bht.scala 200:22]
        btbMeta_40 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_41 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h29 == upIndex) begin // @[bht.scala 200:22]
        btbMeta_41 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_42 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h2a == upIndex) begin // @[bht.scala 200:22]
        btbMeta_42 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_43 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h2b == upIndex) begin // @[bht.scala 200:22]
        btbMeta_43 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_44 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h2c == upIndex) begin // @[bht.scala 200:22]
        btbMeta_44 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_45 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h2d == upIndex) begin // @[bht.scala 200:22]
        btbMeta_45 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_46 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h2e == upIndex) begin // @[bht.scala 200:22]
        btbMeta_46 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_47 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h2f == upIndex) begin // @[bht.scala 200:22]
        btbMeta_47 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_48 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h30 == upIndex) begin // @[bht.scala 200:22]
        btbMeta_48 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_49 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h31 == upIndex) begin // @[bht.scala 200:22]
        btbMeta_49 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_50 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h32 == upIndex) begin // @[bht.scala 200:22]
        btbMeta_50 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_51 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h33 == upIndex) begin // @[bht.scala 200:22]
        btbMeta_51 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_52 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h34 == upIndex) begin // @[bht.scala 200:22]
        btbMeta_52 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_53 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h35 == upIndex) begin // @[bht.scala 200:22]
        btbMeta_53 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_54 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h36 == upIndex) begin // @[bht.scala 200:22]
        btbMeta_54 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_55 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h37 == upIndex) begin // @[bht.scala 200:22]
        btbMeta_55 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_56 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h38 == upIndex) begin // @[bht.scala 200:22]
        btbMeta_56 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_57 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h39 == upIndex) begin // @[bht.scala 200:22]
        btbMeta_57 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_58 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h3a == upIndex) begin // @[bht.scala 200:22]
        btbMeta_58 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_59 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h3b == upIndex) begin // @[bht.scala 200:22]
        btbMeta_59 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_60 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h3c == upIndex) begin // @[bht.scala 200:22]
        btbMeta_60 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_61 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h3d == upIndex) begin // @[bht.scala 200:22]
        btbMeta_61 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_62 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h3e == upIndex) begin // @[bht.scala 200:22]
        btbMeta_62 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_63 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h3f == upIndex) begin // @[bht.scala 200:22]
        btbMeta_63 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_64 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h40 == upIndex) begin // @[bht.scala 200:22]
        btbMeta_64 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_65 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h41 == upIndex) begin // @[bht.scala 200:22]
        btbMeta_65 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_66 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h42 == upIndex) begin // @[bht.scala 200:22]
        btbMeta_66 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_67 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h43 == upIndex) begin // @[bht.scala 200:22]
        btbMeta_67 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_68 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h44 == upIndex) begin // @[bht.scala 200:22]
        btbMeta_68 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_69 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h45 == upIndex) begin // @[bht.scala 200:22]
        btbMeta_69 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_70 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h46 == upIndex) begin // @[bht.scala 200:22]
        btbMeta_70 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_71 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h47 == upIndex) begin // @[bht.scala 200:22]
        btbMeta_71 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_72 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h48 == upIndex) begin // @[bht.scala 200:22]
        btbMeta_72 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_73 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h49 == upIndex) begin // @[bht.scala 200:22]
        btbMeta_73 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_74 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h4a == upIndex) begin // @[bht.scala 200:22]
        btbMeta_74 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_75 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h4b == upIndex) begin // @[bht.scala 200:22]
        btbMeta_75 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_76 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h4c == upIndex) begin // @[bht.scala 200:22]
        btbMeta_76 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_77 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h4d == upIndex) begin // @[bht.scala 200:22]
        btbMeta_77 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_78 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h4e == upIndex) begin // @[bht.scala 200:22]
        btbMeta_78 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_79 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h4f == upIndex) begin // @[bht.scala 200:22]
        btbMeta_79 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_80 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h50 == upIndex) begin // @[bht.scala 200:22]
        btbMeta_80 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_81 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h51 == upIndex) begin // @[bht.scala 200:22]
        btbMeta_81 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_82 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h52 == upIndex) begin // @[bht.scala 200:22]
        btbMeta_82 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_83 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h53 == upIndex) begin // @[bht.scala 200:22]
        btbMeta_83 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_84 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h54 == upIndex) begin // @[bht.scala 200:22]
        btbMeta_84 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_85 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h55 == upIndex) begin // @[bht.scala 200:22]
        btbMeta_85 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_86 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h56 == upIndex) begin // @[bht.scala 200:22]
        btbMeta_86 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_87 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h57 == upIndex) begin // @[bht.scala 200:22]
        btbMeta_87 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_88 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h58 == upIndex) begin // @[bht.scala 200:22]
        btbMeta_88 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_89 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h59 == upIndex) begin // @[bht.scala 200:22]
        btbMeta_89 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_90 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h5a == upIndex) begin // @[bht.scala 200:22]
        btbMeta_90 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_91 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h5b == upIndex) begin // @[bht.scala 200:22]
        btbMeta_91 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_92 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h5c == upIndex) begin // @[bht.scala 200:22]
        btbMeta_92 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_93 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h5d == upIndex) begin // @[bht.scala 200:22]
        btbMeta_93 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_94 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h5e == upIndex) begin // @[bht.scala 200:22]
        btbMeta_94 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_95 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h5f == upIndex) begin // @[bht.scala 200:22]
        btbMeta_95 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_96 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h60 == upIndex) begin // @[bht.scala 200:22]
        btbMeta_96 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_97 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h61 == upIndex) begin // @[bht.scala 200:22]
        btbMeta_97 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_98 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h62 == upIndex) begin // @[bht.scala 200:22]
        btbMeta_98 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_99 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h63 == upIndex) begin // @[bht.scala 200:22]
        btbMeta_99 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_100 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h64 == upIndex) begin // @[bht.scala 200:22]
        btbMeta_100 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_101 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h65 == upIndex) begin // @[bht.scala 200:22]
        btbMeta_101 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_102 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h66 == upIndex) begin // @[bht.scala 200:22]
        btbMeta_102 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_103 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h67 == upIndex) begin // @[bht.scala 200:22]
        btbMeta_103 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_104 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h68 == upIndex) begin // @[bht.scala 200:22]
        btbMeta_104 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_105 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h69 == upIndex) begin // @[bht.scala 200:22]
        btbMeta_105 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_106 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h6a == upIndex) begin // @[bht.scala 200:22]
        btbMeta_106 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_107 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h6b == upIndex) begin // @[bht.scala 200:22]
        btbMeta_107 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_108 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h6c == upIndex) begin // @[bht.scala 200:22]
        btbMeta_108 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_109 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h6d == upIndex) begin // @[bht.scala 200:22]
        btbMeta_109 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_110 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h6e == upIndex) begin // @[bht.scala 200:22]
        btbMeta_110 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_111 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h6f == upIndex) begin // @[bht.scala 200:22]
        btbMeta_111 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_112 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h70 == upIndex) begin // @[bht.scala 200:22]
        btbMeta_112 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_113 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h71 == upIndex) begin // @[bht.scala 200:22]
        btbMeta_113 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_114 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h72 == upIndex) begin // @[bht.scala 200:22]
        btbMeta_114 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_115 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h73 == upIndex) begin // @[bht.scala 200:22]
        btbMeta_115 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_116 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h74 == upIndex) begin // @[bht.scala 200:22]
        btbMeta_116 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_117 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h75 == upIndex) begin // @[bht.scala 200:22]
        btbMeta_117 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_118 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h76 == upIndex) begin // @[bht.scala 200:22]
        btbMeta_118 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_119 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h77 == upIndex) begin // @[bht.scala 200:22]
        btbMeta_119 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_120 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h78 == upIndex) begin // @[bht.scala 200:22]
        btbMeta_120 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_121 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h79 == upIndex) begin // @[bht.scala 200:22]
        btbMeta_121 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_122 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h7a == upIndex) begin // @[bht.scala 200:22]
        btbMeta_122 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_123 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h7b == upIndex) begin // @[bht.scala 200:22]
        btbMeta_123 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_124 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h7c == upIndex) begin // @[bht.scala 200:22]
        btbMeta_124 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_125 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h7d == upIndex) begin // @[bht.scala 200:22]
        btbMeta_125 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_126 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h7e == upIndex) begin // @[bht.scala 200:22]
        btbMeta_126 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    if (reset) begin // @[bht.scala 114:26]
      btbMeta_127 <= 32'h0; // @[bht.scala 114:26]
    end else if (io_fire & (io_takenValid | io_takenValidJalr)) begin // @[bht.scala 196:57]
      if (7'h7f == upIndex) begin // @[bht.scala 200:22]
        btbMeta_127 <= io_nextPC; // @[bht.scala 200:22]
      end
    end
    io_ready_REG <= io_fire; // @[bht.scala 142:48]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ghr = _RAND_0[6:0];
  _RAND_1 = {1{`RANDOM}};
  bht_0 = _RAND_1[6:0];
  _RAND_2 = {1{`RANDOM}};
  bht_1 = _RAND_2[6:0];
  _RAND_3 = {1{`RANDOM}};
  bht_2 = _RAND_3[6:0];
  _RAND_4 = {1{`RANDOM}};
  bht_3 = _RAND_4[6:0];
  _RAND_5 = {1{`RANDOM}};
  bht_4 = _RAND_5[6:0];
  _RAND_6 = {1{`RANDOM}};
  bht_5 = _RAND_6[6:0];
  _RAND_7 = {1{`RANDOM}};
  bht_6 = _RAND_7[6:0];
  _RAND_8 = {1{`RANDOM}};
  bht_7 = _RAND_8[6:0];
  _RAND_9 = {1{`RANDOM}};
  bht_8 = _RAND_9[6:0];
  _RAND_10 = {1{`RANDOM}};
  bht_9 = _RAND_10[6:0];
  _RAND_11 = {1{`RANDOM}};
  bht_10 = _RAND_11[6:0];
  _RAND_12 = {1{`RANDOM}};
  bht_11 = _RAND_12[6:0];
  _RAND_13 = {1{`RANDOM}};
  bht_12 = _RAND_13[6:0];
  _RAND_14 = {1{`RANDOM}};
  bht_13 = _RAND_14[6:0];
  _RAND_15 = {1{`RANDOM}};
  bht_14 = _RAND_15[6:0];
  _RAND_16 = {1{`RANDOM}};
  bht_15 = _RAND_16[6:0];
  _RAND_17 = {1{`RANDOM}};
  bht_16 = _RAND_17[6:0];
  _RAND_18 = {1{`RANDOM}};
  bht_17 = _RAND_18[6:0];
  _RAND_19 = {1{`RANDOM}};
  bht_18 = _RAND_19[6:0];
  _RAND_20 = {1{`RANDOM}};
  bht_19 = _RAND_20[6:0];
  _RAND_21 = {1{`RANDOM}};
  bht_20 = _RAND_21[6:0];
  _RAND_22 = {1{`RANDOM}};
  bht_21 = _RAND_22[6:0];
  _RAND_23 = {1{`RANDOM}};
  bht_22 = _RAND_23[6:0];
  _RAND_24 = {1{`RANDOM}};
  bht_23 = _RAND_24[6:0];
  _RAND_25 = {1{`RANDOM}};
  bht_24 = _RAND_25[6:0];
  _RAND_26 = {1{`RANDOM}};
  bht_25 = _RAND_26[6:0];
  _RAND_27 = {1{`RANDOM}};
  bht_26 = _RAND_27[6:0];
  _RAND_28 = {1{`RANDOM}};
  bht_27 = _RAND_28[6:0];
  _RAND_29 = {1{`RANDOM}};
  bht_28 = _RAND_29[6:0];
  _RAND_30 = {1{`RANDOM}};
  bht_29 = _RAND_30[6:0];
  _RAND_31 = {1{`RANDOM}};
  bht_30 = _RAND_31[6:0];
  _RAND_32 = {1{`RANDOM}};
  bht_31 = _RAND_32[6:0];
  _RAND_33 = {1{`RANDOM}};
  bht_32 = _RAND_33[6:0];
  _RAND_34 = {1{`RANDOM}};
  bht_33 = _RAND_34[6:0];
  _RAND_35 = {1{`RANDOM}};
  bht_34 = _RAND_35[6:0];
  _RAND_36 = {1{`RANDOM}};
  bht_35 = _RAND_36[6:0];
  _RAND_37 = {1{`RANDOM}};
  bht_36 = _RAND_37[6:0];
  _RAND_38 = {1{`RANDOM}};
  bht_37 = _RAND_38[6:0];
  _RAND_39 = {1{`RANDOM}};
  bht_38 = _RAND_39[6:0];
  _RAND_40 = {1{`RANDOM}};
  bht_39 = _RAND_40[6:0];
  _RAND_41 = {1{`RANDOM}};
  bht_40 = _RAND_41[6:0];
  _RAND_42 = {1{`RANDOM}};
  bht_41 = _RAND_42[6:0];
  _RAND_43 = {1{`RANDOM}};
  bht_42 = _RAND_43[6:0];
  _RAND_44 = {1{`RANDOM}};
  bht_43 = _RAND_44[6:0];
  _RAND_45 = {1{`RANDOM}};
  bht_44 = _RAND_45[6:0];
  _RAND_46 = {1{`RANDOM}};
  bht_45 = _RAND_46[6:0];
  _RAND_47 = {1{`RANDOM}};
  bht_46 = _RAND_47[6:0];
  _RAND_48 = {1{`RANDOM}};
  bht_47 = _RAND_48[6:0];
  _RAND_49 = {1{`RANDOM}};
  bht_48 = _RAND_49[6:0];
  _RAND_50 = {1{`RANDOM}};
  bht_49 = _RAND_50[6:0];
  _RAND_51 = {1{`RANDOM}};
  bht_50 = _RAND_51[6:0];
  _RAND_52 = {1{`RANDOM}};
  bht_51 = _RAND_52[6:0];
  _RAND_53 = {1{`RANDOM}};
  bht_52 = _RAND_53[6:0];
  _RAND_54 = {1{`RANDOM}};
  bht_53 = _RAND_54[6:0];
  _RAND_55 = {1{`RANDOM}};
  bht_54 = _RAND_55[6:0];
  _RAND_56 = {1{`RANDOM}};
  bht_55 = _RAND_56[6:0];
  _RAND_57 = {1{`RANDOM}};
  bht_56 = _RAND_57[6:0];
  _RAND_58 = {1{`RANDOM}};
  bht_57 = _RAND_58[6:0];
  _RAND_59 = {1{`RANDOM}};
  bht_58 = _RAND_59[6:0];
  _RAND_60 = {1{`RANDOM}};
  bht_59 = _RAND_60[6:0];
  _RAND_61 = {1{`RANDOM}};
  bht_60 = _RAND_61[6:0];
  _RAND_62 = {1{`RANDOM}};
  bht_61 = _RAND_62[6:0];
  _RAND_63 = {1{`RANDOM}};
  bht_62 = _RAND_63[6:0];
  _RAND_64 = {1{`RANDOM}};
  bht_63 = _RAND_64[6:0];
  _RAND_65 = {1{`RANDOM}};
  bht_64 = _RAND_65[6:0];
  _RAND_66 = {1{`RANDOM}};
  bht_65 = _RAND_66[6:0];
  _RAND_67 = {1{`RANDOM}};
  bht_66 = _RAND_67[6:0];
  _RAND_68 = {1{`RANDOM}};
  bht_67 = _RAND_68[6:0];
  _RAND_69 = {1{`RANDOM}};
  bht_68 = _RAND_69[6:0];
  _RAND_70 = {1{`RANDOM}};
  bht_69 = _RAND_70[6:0];
  _RAND_71 = {1{`RANDOM}};
  bht_70 = _RAND_71[6:0];
  _RAND_72 = {1{`RANDOM}};
  bht_71 = _RAND_72[6:0];
  _RAND_73 = {1{`RANDOM}};
  bht_72 = _RAND_73[6:0];
  _RAND_74 = {1{`RANDOM}};
  bht_73 = _RAND_74[6:0];
  _RAND_75 = {1{`RANDOM}};
  bht_74 = _RAND_75[6:0];
  _RAND_76 = {1{`RANDOM}};
  bht_75 = _RAND_76[6:0];
  _RAND_77 = {1{`RANDOM}};
  bht_76 = _RAND_77[6:0];
  _RAND_78 = {1{`RANDOM}};
  bht_77 = _RAND_78[6:0];
  _RAND_79 = {1{`RANDOM}};
  bht_78 = _RAND_79[6:0];
  _RAND_80 = {1{`RANDOM}};
  bht_79 = _RAND_80[6:0];
  _RAND_81 = {1{`RANDOM}};
  bht_80 = _RAND_81[6:0];
  _RAND_82 = {1{`RANDOM}};
  bht_81 = _RAND_82[6:0];
  _RAND_83 = {1{`RANDOM}};
  bht_82 = _RAND_83[6:0];
  _RAND_84 = {1{`RANDOM}};
  bht_83 = _RAND_84[6:0];
  _RAND_85 = {1{`RANDOM}};
  bht_84 = _RAND_85[6:0];
  _RAND_86 = {1{`RANDOM}};
  bht_85 = _RAND_86[6:0];
  _RAND_87 = {1{`RANDOM}};
  bht_86 = _RAND_87[6:0];
  _RAND_88 = {1{`RANDOM}};
  bht_87 = _RAND_88[6:0];
  _RAND_89 = {1{`RANDOM}};
  bht_88 = _RAND_89[6:0];
  _RAND_90 = {1{`RANDOM}};
  bht_89 = _RAND_90[6:0];
  _RAND_91 = {1{`RANDOM}};
  bht_90 = _RAND_91[6:0];
  _RAND_92 = {1{`RANDOM}};
  bht_91 = _RAND_92[6:0];
  _RAND_93 = {1{`RANDOM}};
  bht_92 = _RAND_93[6:0];
  _RAND_94 = {1{`RANDOM}};
  bht_93 = _RAND_94[6:0];
  _RAND_95 = {1{`RANDOM}};
  bht_94 = _RAND_95[6:0];
  _RAND_96 = {1{`RANDOM}};
  bht_95 = _RAND_96[6:0];
  _RAND_97 = {1{`RANDOM}};
  bht_96 = _RAND_97[6:0];
  _RAND_98 = {1{`RANDOM}};
  bht_97 = _RAND_98[6:0];
  _RAND_99 = {1{`RANDOM}};
  bht_98 = _RAND_99[6:0];
  _RAND_100 = {1{`RANDOM}};
  bht_99 = _RAND_100[6:0];
  _RAND_101 = {1{`RANDOM}};
  bht_100 = _RAND_101[6:0];
  _RAND_102 = {1{`RANDOM}};
  bht_101 = _RAND_102[6:0];
  _RAND_103 = {1{`RANDOM}};
  bht_102 = _RAND_103[6:0];
  _RAND_104 = {1{`RANDOM}};
  bht_103 = _RAND_104[6:0];
  _RAND_105 = {1{`RANDOM}};
  bht_104 = _RAND_105[6:0];
  _RAND_106 = {1{`RANDOM}};
  bht_105 = _RAND_106[6:0];
  _RAND_107 = {1{`RANDOM}};
  bht_106 = _RAND_107[6:0];
  _RAND_108 = {1{`RANDOM}};
  bht_107 = _RAND_108[6:0];
  _RAND_109 = {1{`RANDOM}};
  bht_108 = _RAND_109[6:0];
  _RAND_110 = {1{`RANDOM}};
  bht_109 = _RAND_110[6:0];
  _RAND_111 = {1{`RANDOM}};
  bht_110 = _RAND_111[6:0];
  _RAND_112 = {1{`RANDOM}};
  bht_111 = _RAND_112[6:0];
  _RAND_113 = {1{`RANDOM}};
  bht_112 = _RAND_113[6:0];
  _RAND_114 = {1{`RANDOM}};
  bht_113 = _RAND_114[6:0];
  _RAND_115 = {1{`RANDOM}};
  bht_114 = _RAND_115[6:0];
  _RAND_116 = {1{`RANDOM}};
  bht_115 = _RAND_116[6:0];
  _RAND_117 = {1{`RANDOM}};
  bht_116 = _RAND_117[6:0];
  _RAND_118 = {1{`RANDOM}};
  bht_117 = _RAND_118[6:0];
  _RAND_119 = {1{`RANDOM}};
  bht_118 = _RAND_119[6:0];
  _RAND_120 = {1{`RANDOM}};
  bht_119 = _RAND_120[6:0];
  _RAND_121 = {1{`RANDOM}};
  bht_120 = _RAND_121[6:0];
  _RAND_122 = {1{`RANDOM}};
  bht_121 = _RAND_122[6:0];
  _RAND_123 = {1{`RANDOM}};
  bht_122 = _RAND_123[6:0];
  _RAND_124 = {1{`RANDOM}};
  bht_123 = _RAND_124[6:0];
  _RAND_125 = {1{`RANDOM}};
  bht_124 = _RAND_125[6:0];
  _RAND_126 = {1{`RANDOM}};
  bht_125 = _RAND_126[6:0];
  _RAND_127 = {1{`RANDOM}};
  bht_126 = _RAND_127[6:0];
  _RAND_128 = {1{`RANDOM}};
  bht_127 = _RAND_128[6:0];
  _RAND_129 = {1{`RANDOM}};
  pht_0_0 = _RAND_129[1:0];
  _RAND_130 = {1{`RANDOM}};
  pht_0_1 = _RAND_130[1:0];
  _RAND_131 = {1{`RANDOM}};
  pht_0_2 = _RAND_131[1:0];
  _RAND_132 = {1{`RANDOM}};
  pht_0_3 = _RAND_132[1:0];
  _RAND_133 = {1{`RANDOM}};
  pht_0_4 = _RAND_133[1:0];
  _RAND_134 = {1{`RANDOM}};
  pht_0_5 = _RAND_134[1:0];
  _RAND_135 = {1{`RANDOM}};
  pht_0_6 = _RAND_135[1:0];
  _RAND_136 = {1{`RANDOM}};
  pht_0_7 = _RAND_136[1:0];
  _RAND_137 = {1{`RANDOM}};
  pht_0_8 = _RAND_137[1:0];
  _RAND_138 = {1{`RANDOM}};
  pht_0_9 = _RAND_138[1:0];
  _RAND_139 = {1{`RANDOM}};
  pht_0_10 = _RAND_139[1:0];
  _RAND_140 = {1{`RANDOM}};
  pht_0_11 = _RAND_140[1:0];
  _RAND_141 = {1{`RANDOM}};
  pht_0_12 = _RAND_141[1:0];
  _RAND_142 = {1{`RANDOM}};
  pht_0_13 = _RAND_142[1:0];
  _RAND_143 = {1{`RANDOM}};
  pht_0_14 = _RAND_143[1:0];
  _RAND_144 = {1{`RANDOM}};
  pht_0_15 = _RAND_144[1:0];
  _RAND_145 = {1{`RANDOM}};
  pht_0_16 = _RAND_145[1:0];
  _RAND_146 = {1{`RANDOM}};
  pht_0_17 = _RAND_146[1:0];
  _RAND_147 = {1{`RANDOM}};
  pht_0_18 = _RAND_147[1:0];
  _RAND_148 = {1{`RANDOM}};
  pht_0_19 = _RAND_148[1:0];
  _RAND_149 = {1{`RANDOM}};
  pht_0_20 = _RAND_149[1:0];
  _RAND_150 = {1{`RANDOM}};
  pht_0_21 = _RAND_150[1:0];
  _RAND_151 = {1{`RANDOM}};
  pht_0_22 = _RAND_151[1:0];
  _RAND_152 = {1{`RANDOM}};
  pht_0_23 = _RAND_152[1:0];
  _RAND_153 = {1{`RANDOM}};
  pht_0_24 = _RAND_153[1:0];
  _RAND_154 = {1{`RANDOM}};
  pht_0_25 = _RAND_154[1:0];
  _RAND_155 = {1{`RANDOM}};
  pht_0_26 = _RAND_155[1:0];
  _RAND_156 = {1{`RANDOM}};
  pht_0_27 = _RAND_156[1:0];
  _RAND_157 = {1{`RANDOM}};
  pht_0_28 = _RAND_157[1:0];
  _RAND_158 = {1{`RANDOM}};
  pht_0_29 = _RAND_158[1:0];
  _RAND_159 = {1{`RANDOM}};
  pht_0_30 = _RAND_159[1:0];
  _RAND_160 = {1{`RANDOM}};
  pht_0_31 = _RAND_160[1:0];
  _RAND_161 = {1{`RANDOM}};
  pht_0_32 = _RAND_161[1:0];
  _RAND_162 = {1{`RANDOM}};
  pht_0_33 = _RAND_162[1:0];
  _RAND_163 = {1{`RANDOM}};
  pht_0_34 = _RAND_163[1:0];
  _RAND_164 = {1{`RANDOM}};
  pht_0_35 = _RAND_164[1:0];
  _RAND_165 = {1{`RANDOM}};
  pht_0_36 = _RAND_165[1:0];
  _RAND_166 = {1{`RANDOM}};
  pht_0_37 = _RAND_166[1:0];
  _RAND_167 = {1{`RANDOM}};
  pht_0_38 = _RAND_167[1:0];
  _RAND_168 = {1{`RANDOM}};
  pht_0_39 = _RAND_168[1:0];
  _RAND_169 = {1{`RANDOM}};
  pht_0_40 = _RAND_169[1:0];
  _RAND_170 = {1{`RANDOM}};
  pht_0_41 = _RAND_170[1:0];
  _RAND_171 = {1{`RANDOM}};
  pht_0_42 = _RAND_171[1:0];
  _RAND_172 = {1{`RANDOM}};
  pht_0_43 = _RAND_172[1:0];
  _RAND_173 = {1{`RANDOM}};
  pht_0_44 = _RAND_173[1:0];
  _RAND_174 = {1{`RANDOM}};
  pht_0_45 = _RAND_174[1:0];
  _RAND_175 = {1{`RANDOM}};
  pht_0_46 = _RAND_175[1:0];
  _RAND_176 = {1{`RANDOM}};
  pht_0_47 = _RAND_176[1:0];
  _RAND_177 = {1{`RANDOM}};
  pht_0_48 = _RAND_177[1:0];
  _RAND_178 = {1{`RANDOM}};
  pht_0_49 = _RAND_178[1:0];
  _RAND_179 = {1{`RANDOM}};
  pht_0_50 = _RAND_179[1:0];
  _RAND_180 = {1{`RANDOM}};
  pht_0_51 = _RAND_180[1:0];
  _RAND_181 = {1{`RANDOM}};
  pht_0_52 = _RAND_181[1:0];
  _RAND_182 = {1{`RANDOM}};
  pht_0_53 = _RAND_182[1:0];
  _RAND_183 = {1{`RANDOM}};
  pht_0_54 = _RAND_183[1:0];
  _RAND_184 = {1{`RANDOM}};
  pht_0_55 = _RAND_184[1:0];
  _RAND_185 = {1{`RANDOM}};
  pht_0_56 = _RAND_185[1:0];
  _RAND_186 = {1{`RANDOM}};
  pht_0_57 = _RAND_186[1:0];
  _RAND_187 = {1{`RANDOM}};
  pht_0_58 = _RAND_187[1:0];
  _RAND_188 = {1{`RANDOM}};
  pht_0_59 = _RAND_188[1:0];
  _RAND_189 = {1{`RANDOM}};
  pht_0_60 = _RAND_189[1:0];
  _RAND_190 = {1{`RANDOM}};
  pht_0_61 = _RAND_190[1:0];
  _RAND_191 = {1{`RANDOM}};
  pht_0_62 = _RAND_191[1:0];
  _RAND_192 = {1{`RANDOM}};
  pht_0_63 = _RAND_192[1:0];
  _RAND_193 = {1{`RANDOM}};
  pht_0_64 = _RAND_193[1:0];
  _RAND_194 = {1{`RANDOM}};
  pht_0_65 = _RAND_194[1:0];
  _RAND_195 = {1{`RANDOM}};
  pht_0_66 = _RAND_195[1:0];
  _RAND_196 = {1{`RANDOM}};
  pht_0_67 = _RAND_196[1:0];
  _RAND_197 = {1{`RANDOM}};
  pht_0_68 = _RAND_197[1:0];
  _RAND_198 = {1{`RANDOM}};
  pht_0_69 = _RAND_198[1:0];
  _RAND_199 = {1{`RANDOM}};
  pht_0_70 = _RAND_199[1:0];
  _RAND_200 = {1{`RANDOM}};
  pht_0_71 = _RAND_200[1:0];
  _RAND_201 = {1{`RANDOM}};
  pht_0_72 = _RAND_201[1:0];
  _RAND_202 = {1{`RANDOM}};
  pht_0_73 = _RAND_202[1:0];
  _RAND_203 = {1{`RANDOM}};
  pht_0_74 = _RAND_203[1:0];
  _RAND_204 = {1{`RANDOM}};
  pht_0_75 = _RAND_204[1:0];
  _RAND_205 = {1{`RANDOM}};
  pht_0_76 = _RAND_205[1:0];
  _RAND_206 = {1{`RANDOM}};
  pht_0_77 = _RAND_206[1:0];
  _RAND_207 = {1{`RANDOM}};
  pht_0_78 = _RAND_207[1:0];
  _RAND_208 = {1{`RANDOM}};
  pht_0_79 = _RAND_208[1:0];
  _RAND_209 = {1{`RANDOM}};
  pht_0_80 = _RAND_209[1:0];
  _RAND_210 = {1{`RANDOM}};
  pht_0_81 = _RAND_210[1:0];
  _RAND_211 = {1{`RANDOM}};
  pht_0_82 = _RAND_211[1:0];
  _RAND_212 = {1{`RANDOM}};
  pht_0_83 = _RAND_212[1:0];
  _RAND_213 = {1{`RANDOM}};
  pht_0_84 = _RAND_213[1:0];
  _RAND_214 = {1{`RANDOM}};
  pht_0_85 = _RAND_214[1:0];
  _RAND_215 = {1{`RANDOM}};
  pht_0_86 = _RAND_215[1:0];
  _RAND_216 = {1{`RANDOM}};
  pht_0_87 = _RAND_216[1:0];
  _RAND_217 = {1{`RANDOM}};
  pht_0_88 = _RAND_217[1:0];
  _RAND_218 = {1{`RANDOM}};
  pht_0_89 = _RAND_218[1:0];
  _RAND_219 = {1{`RANDOM}};
  pht_0_90 = _RAND_219[1:0];
  _RAND_220 = {1{`RANDOM}};
  pht_0_91 = _RAND_220[1:0];
  _RAND_221 = {1{`RANDOM}};
  pht_0_92 = _RAND_221[1:0];
  _RAND_222 = {1{`RANDOM}};
  pht_0_93 = _RAND_222[1:0];
  _RAND_223 = {1{`RANDOM}};
  pht_0_94 = _RAND_223[1:0];
  _RAND_224 = {1{`RANDOM}};
  pht_0_95 = _RAND_224[1:0];
  _RAND_225 = {1{`RANDOM}};
  pht_0_96 = _RAND_225[1:0];
  _RAND_226 = {1{`RANDOM}};
  pht_0_97 = _RAND_226[1:0];
  _RAND_227 = {1{`RANDOM}};
  pht_0_98 = _RAND_227[1:0];
  _RAND_228 = {1{`RANDOM}};
  pht_0_99 = _RAND_228[1:0];
  _RAND_229 = {1{`RANDOM}};
  pht_0_100 = _RAND_229[1:0];
  _RAND_230 = {1{`RANDOM}};
  pht_0_101 = _RAND_230[1:0];
  _RAND_231 = {1{`RANDOM}};
  pht_0_102 = _RAND_231[1:0];
  _RAND_232 = {1{`RANDOM}};
  pht_0_103 = _RAND_232[1:0];
  _RAND_233 = {1{`RANDOM}};
  pht_0_104 = _RAND_233[1:0];
  _RAND_234 = {1{`RANDOM}};
  pht_0_105 = _RAND_234[1:0];
  _RAND_235 = {1{`RANDOM}};
  pht_0_106 = _RAND_235[1:0];
  _RAND_236 = {1{`RANDOM}};
  pht_0_107 = _RAND_236[1:0];
  _RAND_237 = {1{`RANDOM}};
  pht_0_108 = _RAND_237[1:0];
  _RAND_238 = {1{`RANDOM}};
  pht_0_109 = _RAND_238[1:0];
  _RAND_239 = {1{`RANDOM}};
  pht_0_110 = _RAND_239[1:0];
  _RAND_240 = {1{`RANDOM}};
  pht_0_111 = _RAND_240[1:0];
  _RAND_241 = {1{`RANDOM}};
  pht_0_112 = _RAND_241[1:0];
  _RAND_242 = {1{`RANDOM}};
  pht_0_113 = _RAND_242[1:0];
  _RAND_243 = {1{`RANDOM}};
  pht_0_114 = _RAND_243[1:0];
  _RAND_244 = {1{`RANDOM}};
  pht_0_115 = _RAND_244[1:0];
  _RAND_245 = {1{`RANDOM}};
  pht_0_116 = _RAND_245[1:0];
  _RAND_246 = {1{`RANDOM}};
  pht_0_117 = _RAND_246[1:0];
  _RAND_247 = {1{`RANDOM}};
  pht_0_118 = _RAND_247[1:0];
  _RAND_248 = {1{`RANDOM}};
  pht_0_119 = _RAND_248[1:0];
  _RAND_249 = {1{`RANDOM}};
  pht_0_120 = _RAND_249[1:0];
  _RAND_250 = {1{`RANDOM}};
  pht_0_121 = _RAND_250[1:0];
  _RAND_251 = {1{`RANDOM}};
  pht_0_122 = _RAND_251[1:0];
  _RAND_252 = {1{`RANDOM}};
  pht_0_123 = _RAND_252[1:0];
  _RAND_253 = {1{`RANDOM}};
  pht_0_124 = _RAND_253[1:0];
  _RAND_254 = {1{`RANDOM}};
  pht_0_125 = _RAND_254[1:0];
  _RAND_255 = {1{`RANDOM}};
  pht_0_126 = _RAND_255[1:0];
  _RAND_256 = {1{`RANDOM}};
  pht_0_127 = _RAND_256[1:0];
  _RAND_257 = {1{`RANDOM}};
  pht_1_0 = _RAND_257[1:0];
  _RAND_258 = {1{`RANDOM}};
  pht_1_1 = _RAND_258[1:0];
  _RAND_259 = {1{`RANDOM}};
  pht_1_2 = _RAND_259[1:0];
  _RAND_260 = {1{`RANDOM}};
  pht_1_3 = _RAND_260[1:0];
  _RAND_261 = {1{`RANDOM}};
  pht_1_4 = _RAND_261[1:0];
  _RAND_262 = {1{`RANDOM}};
  pht_1_5 = _RAND_262[1:0];
  _RAND_263 = {1{`RANDOM}};
  pht_1_6 = _RAND_263[1:0];
  _RAND_264 = {1{`RANDOM}};
  pht_1_7 = _RAND_264[1:0];
  _RAND_265 = {1{`RANDOM}};
  pht_1_8 = _RAND_265[1:0];
  _RAND_266 = {1{`RANDOM}};
  pht_1_9 = _RAND_266[1:0];
  _RAND_267 = {1{`RANDOM}};
  pht_1_10 = _RAND_267[1:0];
  _RAND_268 = {1{`RANDOM}};
  pht_1_11 = _RAND_268[1:0];
  _RAND_269 = {1{`RANDOM}};
  pht_1_12 = _RAND_269[1:0];
  _RAND_270 = {1{`RANDOM}};
  pht_1_13 = _RAND_270[1:0];
  _RAND_271 = {1{`RANDOM}};
  pht_1_14 = _RAND_271[1:0];
  _RAND_272 = {1{`RANDOM}};
  pht_1_15 = _RAND_272[1:0];
  _RAND_273 = {1{`RANDOM}};
  pht_1_16 = _RAND_273[1:0];
  _RAND_274 = {1{`RANDOM}};
  pht_1_17 = _RAND_274[1:0];
  _RAND_275 = {1{`RANDOM}};
  pht_1_18 = _RAND_275[1:0];
  _RAND_276 = {1{`RANDOM}};
  pht_1_19 = _RAND_276[1:0];
  _RAND_277 = {1{`RANDOM}};
  pht_1_20 = _RAND_277[1:0];
  _RAND_278 = {1{`RANDOM}};
  pht_1_21 = _RAND_278[1:0];
  _RAND_279 = {1{`RANDOM}};
  pht_1_22 = _RAND_279[1:0];
  _RAND_280 = {1{`RANDOM}};
  pht_1_23 = _RAND_280[1:0];
  _RAND_281 = {1{`RANDOM}};
  pht_1_24 = _RAND_281[1:0];
  _RAND_282 = {1{`RANDOM}};
  pht_1_25 = _RAND_282[1:0];
  _RAND_283 = {1{`RANDOM}};
  pht_1_26 = _RAND_283[1:0];
  _RAND_284 = {1{`RANDOM}};
  pht_1_27 = _RAND_284[1:0];
  _RAND_285 = {1{`RANDOM}};
  pht_1_28 = _RAND_285[1:0];
  _RAND_286 = {1{`RANDOM}};
  pht_1_29 = _RAND_286[1:0];
  _RAND_287 = {1{`RANDOM}};
  pht_1_30 = _RAND_287[1:0];
  _RAND_288 = {1{`RANDOM}};
  pht_1_31 = _RAND_288[1:0];
  _RAND_289 = {1{`RANDOM}};
  pht_1_32 = _RAND_289[1:0];
  _RAND_290 = {1{`RANDOM}};
  pht_1_33 = _RAND_290[1:0];
  _RAND_291 = {1{`RANDOM}};
  pht_1_34 = _RAND_291[1:0];
  _RAND_292 = {1{`RANDOM}};
  pht_1_35 = _RAND_292[1:0];
  _RAND_293 = {1{`RANDOM}};
  pht_1_36 = _RAND_293[1:0];
  _RAND_294 = {1{`RANDOM}};
  pht_1_37 = _RAND_294[1:0];
  _RAND_295 = {1{`RANDOM}};
  pht_1_38 = _RAND_295[1:0];
  _RAND_296 = {1{`RANDOM}};
  pht_1_39 = _RAND_296[1:0];
  _RAND_297 = {1{`RANDOM}};
  pht_1_40 = _RAND_297[1:0];
  _RAND_298 = {1{`RANDOM}};
  pht_1_41 = _RAND_298[1:0];
  _RAND_299 = {1{`RANDOM}};
  pht_1_42 = _RAND_299[1:0];
  _RAND_300 = {1{`RANDOM}};
  pht_1_43 = _RAND_300[1:0];
  _RAND_301 = {1{`RANDOM}};
  pht_1_44 = _RAND_301[1:0];
  _RAND_302 = {1{`RANDOM}};
  pht_1_45 = _RAND_302[1:0];
  _RAND_303 = {1{`RANDOM}};
  pht_1_46 = _RAND_303[1:0];
  _RAND_304 = {1{`RANDOM}};
  pht_1_47 = _RAND_304[1:0];
  _RAND_305 = {1{`RANDOM}};
  pht_1_48 = _RAND_305[1:0];
  _RAND_306 = {1{`RANDOM}};
  pht_1_49 = _RAND_306[1:0];
  _RAND_307 = {1{`RANDOM}};
  pht_1_50 = _RAND_307[1:0];
  _RAND_308 = {1{`RANDOM}};
  pht_1_51 = _RAND_308[1:0];
  _RAND_309 = {1{`RANDOM}};
  pht_1_52 = _RAND_309[1:0];
  _RAND_310 = {1{`RANDOM}};
  pht_1_53 = _RAND_310[1:0];
  _RAND_311 = {1{`RANDOM}};
  pht_1_54 = _RAND_311[1:0];
  _RAND_312 = {1{`RANDOM}};
  pht_1_55 = _RAND_312[1:0];
  _RAND_313 = {1{`RANDOM}};
  pht_1_56 = _RAND_313[1:0];
  _RAND_314 = {1{`RANDOM}};
  pht_1_57 = _RAND_314[1:0];
  _RAND_315 = {1{`RANDOM}};
  pht_1_58 = _RAND_315[1:0];
  _RAND_316 = {1{`RANDOM}};
  pht_1_59 = _RAND_316[1:0];
  _RAND_317 = {1{`RANDOM}};
  pht_1_60 = _RAND_317[1:0];
  _RAND_318 = {1{`RANDOM}};
  pht_1_61 = _RAND_318[1:0];
  _RAND_319 = {1{`RANDOM}};
  pht_1_62 = _RAND_319[1:0];
  _RAND_320 = {1{`RANDOM}};
  pht_1_63 = _RAND_320[1:0];
  _RAND_321 = {1{`RANDOM}};
  pht_1_64 = _RAND_321[1:0];
  _RAND_322 = {1{`RANDOM}};
  pht_1_65 = _RAND_322[1:0];
  _RAND_323 = {1{`RANDOM}};
  pht_1_66 = _RAND_323[1:0];
  _RAND_324 = {1{`RANDOM}};
  pht_1_67 = _RAND_324[1:0];
  _RAND_325 = {1{`RANDOM}};
  pht_1_68 = _RAND_325[1:0];
  _RAND_326 = {1{`RANDOM}};
  pht_1_69 = _RAND_326[1:0];
  _RAND_327 = {1{`RANDOM}};
  pht_1_70 = _RAND_327[1:0];
  _RAND_328 = {1{`RANDOM}};
  pht_1_71 = _RAND_328[1:0];
  _RAND_329 = {1{`RANDOM}};
  pht_1_72 = _RAND_329[1:0];
  _RAND_330 = {1{`RANDOM}};
  pht_1_73 = _RAND_330[1:0];
  _RAND_331 = {1{`RANDOM}};
  pht_1_74 = _RAND_331[1:0];
  _RAND_332 = {1{`RANDOM}};
  pht_1_75 = _RAND_332[1:0];
  _RAND_333 = {1{`RANDOM}};
  pht_1_76 = _RAND_333[1:0];
  _RAND_334 = {1{`RANDOM}};
  pht_1_77 = _RAND_334[1:0];
  _RAND_335 = {1{`RANDOM}};
  pht_1_78 = _RAND_335[1:0];
  _RAND_336 = {1{`RANDOM}};
  pht_1_79 = _RAND_336[1:0];
  _RAND_337 = {1{`RANDOM}};
  pht_1_80 = _RAND_337[1:0];
  _RAND_338 = {1{`RANDOM}};
  pht_1_81 = _RAND_338[1:0];
  _RAND_339 = {1{`RANDOM}};
  pht_1_82 = _RAND_339[1:0];
  _RAND_340 = {1{`RANDOM}};
  pht_1_83 = _RAND_340[1:0];
  _RAND_341 = {1{`RANDOM}};
  pht_1_84 = _RAND_341[1:0];
  _RAND_342 = {1{`RANDOM}};
  pht_1_85 = _RAND_342[1:0];
  _RAND_343 = {1{`RANDOM}};
  pht_1_86 = _RAND_343[1:0];
  _RAND_344 = {1{`RANDOM}};
  pht_1_87 = _RAND_344[1:0];
  _RAND_345 = {1{`RANDOM}};
  pht_1_88 = _RAND_345[1:0];
  _RAND_346 = {1{`RANDOM}};
  pht_1_89 = _RAND_346[1:0];
  _RAND_347 = {1{`RANDOM}};
  pht_1_90 = _RAND_347[1:0];
  _RAND_348 = {1{`RANDOM}};
  pht_1_91 = _RAND_348[1:0];
  _RAND_349 = {1{`RANDOM}};
  pht_1_92 = _RAND_349[1:0];
  _RAND_350 = {1{`RANDOM}};
  pht_1_93 = _RAND_350[1:0];
  _RAND_351 = {1{`RANDOM}};
  pht_1_94 = _RAND_351[1:0];
  _RAND_352 = {1{`RANDOM}};
  pht_1_95 = _RAND_352[1:0];
  _RAND_353 = {1{`RANDOM}};
  pht_1_96 = _RAND_353[1:0];
  _RAND_354 = {1{`RANDOM}};
  pht_1_97 = _RAND_354[1:0];
  _RAND_355 = {1{`RANDOM}};
  pht_1_98 = _RAND_355[1:0];
  _RAND_356 = {1{`RANDOM}};
  pht_1_99 = _RAND_356[1:0];
  _RAND_357 = {1{`RANDOM}};
  pht_1_100 = _RAND_357[1:0];
  _RAND_358 = {1{`RANDOM}};
  pht_1_101 = _RAND_358[1:0];
  _RAND_359 = {1{`RANDOM}};
  pht_1_102 = _RAND_359[1:0];
  _RAND_360 = {1{`RANDOM}};
  pht_1_103 = _RAND_360[1:0];
  _RAND_361 = {1{`RANDOM}};
  pht_1_104 = _RAND_361[1:0];
  _RAND_362 = {1{`RANDOM}};
  pht_1_105 = _RAND_362[1:0];
  _RAND_363 = {1{`RANDOM}};
  pht_1_106 = _RAND_363[1:0];
  _RAND_364 = {1{`RANDOM}};
  pht_1_107 = _RAND_364[1:0];
  _RAND_365 = {1{`RANDOM}};
  pht_1_108 = _RAND_365[1:0];
  _RAND_366 = {1{`RANDOM}};
  pht_1_109 = _RAND_366[1:0];
  _RAND_367 = {1{`RANDOM}};
  pht_1_110 = _RAND_367[1:0];
  _RAND_368 = {1{`RANDOM}};
  pht_1_111 = _RAND_368[1:0];
  _RAND_369 = {1{`RANDOM}};
  pht_1_112 = _RAND_369[1:0];
  _RAND_370 = {1{`RANDOM}};
  pht_1_113 = _RAND_370[1:0];
  _RAND_371 = {1{`RANDOM}};
  pht_1_114 = _RAND_371[1:0];
  _RAND_372 = {1{`RANDOM}};
  pht_1_115 = _RAND_372[1:0];
  _RAND_373 = {1{`RANDOM}};
  pht_1_116 = _RAND_373[1:0];
  _RAND_374 = {1{`RANDOM}};
  pht_1_117 = _RAND_374[1:0];
  _RAND_375 = {1{`RANDOM}};
  pht_1_118 = _RAND_375[1:0];
  _RAND_376 = {1{`RANDOM}};
  pht_1_119 = _RAND_376[1:0];
  _RAND_377 = {1{`RANDOM}};
  pht_1_120 = _RAND_377[1:0];
  _RAND_378 = {1{`RANDOM}};
  pht_1_121 = _RAND_378[1:0];
  _RAND_379 = {1{`RANDOM}};
  pht_1_122 = _RAND_379[1:0];
  _RAND_380 = {1{`RANDOM}};
  pht_1_123 = _RAND_380[1:0];
  _RAND_381 = {1{`RANDOM}};
  pht_1_124 = _RAND_381[1:0];
  _RAND_382 = {1{`RANDOM}};
  pht_1_125 = _RAND_382[1:0];
  _RAND_383 = {1{`RANDOM}};
  pht_1_126 = _RAND_383[1:0];
  _RAND_384 = {1{`RANDOM}};
  pht_1_127 = _RAND_384[1:0];
  _RAND_385 = {1{`RANDOM}};
  pht_2_0 = _RAND_385[1:0];
  _RAND_386 = {1{`RANDOM}};
  pht_2_1 = _RAND_386[1:0];
  _RAND_387 = {1{`RANDOM}};
  pht_2_2 = _RAND_387[1:0];
  _RAND_388 = {1{`RANDOM}};
  pht_2_3 = _RAND_388[1:0];
  _RAND_389 = {1{`RANDOM}};
  pht_2_4 = _RAND_389[1:0];
  _RAND_390 = {1{`RANDOM}};
  pht_2_5 = _RAND_390[1:0];
  _RAND_391 = {1{`RANDOM}};
  pht_2_6 = _RAND_391[1:0];
  _RAND_392 = {1{`RANDOM}};
  pht_2_7 = _RAND_392[1:0];
  _RAND_393 = {1{`RANDOM}};
  pht_2_8 = _RAND_393[1:0];
  _RAND_394 = {1{`RANDOM}};
  pht_2_9 = _RAND_394[1:0];
  _RAND_395 = {1{`RANDOM}};
  pht_2_10 = _RAND_395[1:0];
  _RAND_396 = {1{`RANDOM}};
  pht_2_11 = _RAND_396[1:0];
  _RAND_397 = {1{`RANDOM}};
  pht_2_12 = _RAND_397[1:0];
  _RAND_398 = {1{`RANDOM}};
  pht_2_13 = _RAND_398[1:0];
  _RAND_399 = {1{`RANDOM}};
  pht_2_14 = _RAND_399[1:0];
  _RAND_400 = {1{`RANDOM}};
  pht_2_15 = _RAND_400[1:0];
  _RAND_401 = {1{`RANDOM}};
  pht_2_16 = _RAND_401[1:0];
  _RAND_402 = {1{`RANDOM}};
  pht_2_17 = _RAND_402[1:0];
  _RAND_403 = {1{`RANDOM}};
  pht_2_18 = _RAND_403[1:0];
  _RAND_404 = {1{`RANDOM}};
  pht_2_19 = _RAND_404[1:0];
  _RAND_405 = {1{`RANDOM}};
  pht_2_20 = _RAND_405[1:0];
  _RAND_406 = {1{`RANDOM}};
  pht_2_21 = _RAND_406[1:0];
  _RAND_407 = {1{`RANDOM}};
  pht_2_22 = _RAND_407[1:0];
  _RAND_408 = {1{`RANDOM}};
  pht_2_23 = _RAND_408[1:0];
  _RAND_409 = {1{`RANDOM}};
  pht_2_24 = _RAND_409[1:0];
  _RAND_410 = {1{`RANDOM}};
  pht_2_25 = _RAND_410[1:0];
  _RAND_411 = {1{`RANDOM}};
  pht_2_26 = _RAND_411[1:0];
  _RAND_412 = {1{`RANDOM}};
  pht_2_27 = _RAND_412[1:0];
  _RAND_413 = {1{`RANDOM}};
  pht_2_28 = _RAND_413[1:0];
  _RAND_414 = {1{`RANDOM}};
  pht_2_29 = _RAND_414[1:0];
  _RAND_415 = {1{`RANDOM}};
  pht_2_30 = _RAND_415[1:0];
  _RAND_416 = {1{`RANDOM}};
  pht_2_31 = _RAND_416[1:0];
  _RAND_417 = {1{`RANDOM}};
  pht_2_32 = _RAND_417[1:0];
  _RAND_418 = {1{`RANDOM}};
  pht_2_33 = _RAND_418[1:0];
  _RAND_419 = {1{`RANDOM}};
  pht_2_34 = _RAND_419[1:0];
  _RAND_420 = {1{`RANDOM}};
  pht_2_35 = _RAND_420[1:0];
  _RAND_421 = {1{`RANDOM}};
  pht_2_36 = _RAND_421[1:0];
  _RAND_422 = {1{`RANDOM}};
  pht_2_37 = _RAND_422[1:0];
  _RAND_423 = {1{`RANDOM}};
  pht_2_38 = _RAND_423[1:0];
  _RAND_424 = {1{`RANDOM}};
  pht_2_39 = _RAND_424[1:0];
  _RAND_425 = {1{`RANDOM}};
  pht_2_40 = _RAND_425[1:0];
  _RAND_426 = {1{`RANDOM}};
  pht_2_41 = _RAND_426[1:0];
  _RAND_427 = {1{`RANDOM}};
  pht_2_42 = _RAND_427[1:0];
  _RAND_428 = {1{`RANDOM}};
  pht_2_43 = _RAND_428[1:0];
  _RAND_429 = {1{`RANDOM}};
  pht_2_44 = _RAND_429[1:0];
  _RAND_430 = {1{`RANDOM}};
  pht_2_45 = _RAND_430[1:0];
  _RAND_431 = {1{`RANDOM}};
  pht_2_46 = _RAND_431[1:0];
  _RAND_432 = {1{`RANDOM}};
  pht_2_47 = _RAND_432[1:0];
  _RAND_433 = {1{`RANDOM}};
  pht_2_48 = _RAND_433[1:0];
  _RAND_434 = {1{`RANDOM}};
  pht_2_49 = _RAND_434[1:0];
  _RAND_435 = {1{`RANDOM}};
  pht_2_50 = _RAND_435[1:0];
  _RAND_436 = {1{`RANDOM}};
  pht_2_51 = _RAND_436[1:0];
  _RAND_437 = {1{`RANDOM}};
  pht_2_52 = _RAND_437[1:0];
  _RAND_438 = {1{`RANDOM}};
  pht_2_53 = _RAND_438[1:0];
  _RAND_439 = {1{`RANDOM}};
  pht_2_54 = _RAND_439[1:0];
  _RAND_440 = {1{`RANDOM}};
  pht_2_55 = _RAND_440[1:0];
  _RAND_441 = {1{`RANDOM}};
  pht_2_56 = _RAND_441[1:0];
  _RAND_442 = {1{`RANDOM}};
  pht_2_57 = _RAND_442[1:0];
  _RAND_443 = {1{`RANDOM}};
  pht_2_58 = _RAND_443[1:0];
  _RAND_444 = {1{`RANDOM}};
  pht_2_59 = _RAND_444[1:0];
  _RAND_445 = {1{`RANDOM}};
  pht_2_60 = _RAND_445[1:0];
  _RAND_446 = {1{`RANDOM}};
  pht_2_61 = _RAND_446[1:0];
  _RAND_447 = {1{`RANDOM}};
  pht_2_62 = _RAND_447[1:0];
  _RAND_448 = {1{`RANDOM}};
  pht_2_63 = _RAND_448[1:0];
  _RAND_449 = {1{`RANDOM}};
  pht_2_64 = _RAND_449[1:0];
  _RAND_450 = {1{`RANDOM}};
  pht_2_65 = _RAND_450[1:0];
  _RAND_451 = {1{`RANDOM}};
  pht_2_66 = _RAND_451[1:0];
  _RAND_452 = {1{`RANDOM}};
  pht_2_67 = _RAND_452[1:0];
  _RAND_453 = {1{`RANDOM}};
  pht_2_68 = _RAND_453[1:0];
  _RAND_454 = {1{`RANDOM}};
  pht_2_69 = _RAND_454[1:0];
  _RAND_455 = {1{`RANDOM}};
  pht_2_70 = _RAND_455[1:0];
  _RAND_456 = {1{`RANDOM}};
  pht_2_71 = _RAND_456[1:0];
  _RAND_457 = {1{`RANDOM}};
  pht_2_72 = _RAND_457[1:0];
  _RAND_458 = {1{`RANDOM}};
  pht_2_73 = _RAND_458[1:0];
  _RAND_459 = {1{`RANDOM}};
  pht_2_74 = _RAND_459[1:0];
  _RAND_460 = {1{`RANDOM}};
  pht_2_75 = _RAND_460[1:0];
  _RAND_461 = {1{`RANDOM}};
  pht_2_76 = _RAND_461[1:0];
  _RAND_462 = {1{`RANDOM}};
  pht_2_77 = _RAND_462[1:0];
  _RAND_463 = {1{`RANDOM}};
  pht_2_78 = _RAND_463[1:0];
  _RAND_464 = {1{`RANDOM}};
  pht_2_79 = _RAND_464[1:0];
  _RAND_465 = {1{`RANDOM}};
  pht_2_80 = _RAND_465[1:0];
  _RAND_466 = {1{`RANDOM}};
  pht_2_81 = _RAND_466[1:0];
  _RAND_467 = {1{`RANDOM}};
  pht_2_82 = _RAND_467[1:0];
  _RAND_468 = {1{`RANDOM}};
  pht_2_83 = _RAND_468[1:0];
  _RAND_469 = {1{`RANDOM}};
  pht_2_84 = _RAND_469[1:0];
  _RAND_470 = {1{`RANDOM}};
  pht_2_85 = _RAND_470[1:0];
  _RAND_471 = {1{`RANDOM}};
  pht_2_86 = _RAND_471[1:0];
  _RAND_472 = {1{`RANDOM}};
  pht_2_87 = _RAND_472[1:0];
  _RAND_473 = {1{`RANDOM}};
  pht_2_88 = _RAND_473[1:0];
  _RAND_474 = {1{`RANDOM}};
  pht_2_89 = _RAND_474[1:0];
  _RAND_475 = {1{`RANDOM}};
  pht_2_90 = _RAND_475[1:0];
  _RAND_476 = {1{`RANDOM}};
  pht_2_91 = _RAND_476[1:0];
  _RAND_477 = {1{`RANDOM}};
  pht_2_92 = _RAND_477[1:0];
  _RAND_478 = {1{`RANDOM}};
  pht_2_93 = _RAND_478[1:0];
  _RAND_479 = {1{`RANDOM}};
  pht_2_94 = _RAND_479[1:0];
  _RAND_480 = {1{`RANDOM}};
  pht_2_95 = _RAND_480[1:0];
  _RAND_481 = {1{`RANDOM}};
  pht_2_96 = _RAND_481[1:0];
  _RAND_482 = {1{`RANDOM}};
  pht_2_97 = _RAND_482[1:0];
  _RAND_483 = {1{`RANDOM}};
  pht_2_98 = _RAND_483[1:0];
  _RAND_484 = {1{`RANDOM}};
  pht_2_99 = _RAND_484[1:0];
  _RAND_485 = {1{`RANDOM}};
  pht_2_100 = _RAND_485[1:0];
  _RAND_486 = {1{`RANDOM}};
  pht_2_101 = _RAND_486[1:0];
  _RAND_487 = {1{`RANDOM}};
  pht_2_102 = _RAND_487[1:0];
  _RAND_488 = {1{`RANDOM}};
  pht_2_103 = _RAND_488[1:0];
  _RAND_489 = {1{`RANDOM}};
  pht_2_104 = _RAND_489[1:0];
  _RAND_490 = {1{`RANDOM}};
  pht_2_105 = _RAND_490[1:0];
  _RAND_491 = {1{`RANDOM}};
  pht_2_106 = _RAND_491[1:0];
  _RAND_492 = {1{`RANDOM}};
  pht_2_107 = _RAND_492[1:0];
  _RAND_493 = {1{`RANDOM}};
  pht_2_108 = _RAND_493[1:0];
  _RAND_494 = {1{`RANDOM}};
  pht_2_109 = _RAND_494[1:0];
  _RAND_495 = {1{`RANDOM}};
  pht_2_110 = _RAND_495[1:0];
  _RAND_496 = {1{`RANDOM}};
  pht_2_111 = _RAND_496[1:0];
  _RAND_497 = {1{`RANDOM}};
  pht_2_112 = _RAND_497[1:0];
  _RAND_498 = {1{`RANDOM}};
  pht_2_113 = _RAND_498[1:0];
  _RAND_499 = {1{`RANDOM}};
  pht_2_114 = _RAND_499[1:0];
  _RAND_500 = {1{`RANDOM}};
  pht_2_115 = _RAND_500[1:0];
  _RAND_501 = {1{`RANDOM}};
  pht_2_116 = _RAND_501[1:0];
  _RAND_502 = {1{`RANDOM}};
  pht_2_117 = _RAND_502[1:0];
  _RAND_503 = {1{`RANDOM}};
  pht_2_118 = _RAND_503[1:0];
  _RAND_504 = {1{`RANDOM}};
  pht_2_119 = _RAND_504[1:0];
  _RAND_505 = {1{`RANDOM}};
  pht_2_120 = _RAND_505[1:0];
  _RAND_506 = {1{`RANDOM}};
  pht_2_121 = _RAND_506[1:0];
  _RAND_507 = {1{`RANDOM}};
  pht_2_122 = _RAND_507[1:0];
  _RAND_508 = {1{`RANDOM}};
  pht_2_123 = _RAND_508[1:0];
  _RAND_509 = {1{`RANDOM}};
  pht_2_124 = _RAND_509[1:0];
  _RAND_510 = {1{`RANDOM}};
  pht_2_125 = _RAND_510[1:0];
  _RAND_511 = {1{`RANDOM}};
  pht_2_126 = _RAND_511[1:0];
  _RAND_512 = {1{`RANDOM}};
  pht_2_127 = _RAND_512[1:0];
  _RAND_513 = {1{`RANDOM}};
  btbV_0 = _RAND_513[0:0];
  _RAND_514 = {1{`RANDOM}};
  btbV_1 = _RAND_514[0:0];
  _RAND_515 = {1{`RANDOM}};
  btbV_2 = _RAND_515[0:0];
  _RAND_516 = {1{`RANDOM}};
  btbV_3 = _RAND_516[0:0];
  _RAND_517 = {1{`RANDOM}};
  btbV_4 = _RAND_517[0:0];
  _RAND_518 = {1{`RANDOM}};
  btbV_5 = _RAND_518[0:0];
  _RAND_519 = {1{`RANDOM}};
  btbV_6 = _RAND_519[0:0];
  _RAND_520 = {1{`RANDOM}};
  btbV_7 = _RAND_520[0:0];
  _RAND_521 = {1{`RANDOM}};
  btbV_8 = _RAND_521[0:0];
  _RAND_522 = {1{`RANDOM}};
  btbV_9 = _RAND_522[0:0];
  _RAND_523 = {1{`RANDOM}};
  btbV_10 = _RAND_523[0:0];
  _RAND_524 = {1{`RANDOM}};
  btbV_11 = _RAND_524[0:0];
  _RAND_525 = {1{`RANDOM}};
  btbV_12 = _RAND_525[0:0];
  _RAND_526 = {1{`RANDOM}};
  btbV_13 = _RAND_526[0:0];
  _RAND_527 = {1{`RANDOM}};
  btbV_14 = _RAND_527[0:0];
  _RAND_528 = {1{`RANDOM}};
  btbV_15 = _RAND_528[0:0];
  _RAND_529 = {1{`RANDOM}};
  btbV_16 = _RAND_529[0:0];
  _RAND_530 = {1{`RANDOM}};
  btbV_17 = _RAND_530[0:0];
  _RAND_531 = {1{`RANDOM}};
  btbV_18 = _RAND_531[0:0];
  _RAND_532 = {1{`RANDOM}};
  btbV_19 = _RAND_532[0:0];
  _RAND_533 = {1{`RANDOM}};
  btbV_20 = _RAND_533[0:0];
  _RAND_534 = {1{`RANDOM}};
  btbV_21 = _RAND_534[0:0];
  _RAND_535 = {1{`RANDOM}};
  btbV_22 = _RAND_535[0:0];
  _RAND_536 = {1{`RANDOM}};
  btbV_23 = _RAND_536[0:0];
  _RAND_537 = {1{`RANDOM}};
  btbV_24 = _RAND_537[0:0];
  _RAND_538 = {1{`RANDOM}};
  btbV_25 = _RAND_538[0:0];
  _RAND_539 = {1{`RANDOM}};
  btbV_26 = _RAND_539[0:0];
  _RAND_540 = {1{`RANDOM}};
  btbV_27 = _RAND_540[0:0];
  _RAND_541 = {1{`RANDOM}};
  btbV_28 = _RAND_541[0:0];
  _RAND_542 = {1{`RANDOM}};
  btbV_29 = _RAND_542[0:0];
  _RAND_543 = {1{`RANDOM}};
  btbV_30 = _RAND_543[0:0];
  _RAND_544 = {1{`RANDOM}};
  btbV_31 = _RAND_544[0:0];
  _RAND_545 = {1{`RANDOM}};
  btbV_32 = _RAND_545[0:0];
  _RAND_546 = {1{`RANDOM}};
  btbV_33 = _RAND_546[0:0];
  _RAND_547 = {1{`RANDOM}};
  btbV_34 = _RAND_547[0:0];
  _RAND_548 = {1{`RANDOM}};
  btbV_35 = _RAND_548[0:0];
  _RAND_549 = {1{`RANDOM}};
  btbV_36 = _RAND_549[0:0];
  _RAND_550 = {1{`RANDOM}};
  btbV_37 = _RAND_550[0:0];
  _RAND_551 = {1{`RANDOM}};
  btbV_38 = _RAND_551[0:0];
  _RAND_552 = {1{`RANDOM}};
  btbV_39 = _RAND_552[0:0];
  _RAND_553 = {1{`RANDOM}};
  btbV_40 = _RAND_553[0:0];
  _RAND_554 = {1{`RANDOM}};
  btbV_41 = _RAND_554[0:0];
  _RAND_555 = {1{`RANDOM}};
  btbV_42 = _RAND_555[0:0];
  _RAND_556 = {1{`RANDOM}};
  btbV_43 = _RAND_556[0:0];
  _RAND_557 = {1{`RANDOM}};
  btbV_44 = _RAND_557[0:0];
  _RAND_558 = {1{`RANDOM}};
  btbV_45 = _RAND_558[0:0];
  _RAND_559 = {1{`RANDOM}};
  btbV_46 = _RAND_559[0:0];
  _RAND_560 = {1{`RANDOM}};
  btbV_47 = _RAND_560[0:0];
  _RAND_561 = {1{`RANDOM}};
  btbV_48 = _RAND_561[0:0];
  _RAND_562 = {1{`RANDOM}};
  btbV_49 = _RAND_562[0:0];
  _RAND_563 = {1{`RANDOM}};
  btbV_50 = _RAND_563[0:0];
  _RAND_564 = {1{`RANDOM}};
  btbV_51 = _RAND_564[0:0];
  _RAND_565 = {1{`RANDOM}};
  btbV_52 = _RAND_565[0:0];
  _RAND_566 = {1{`RANDOM}};
  btbV_53 = _RAND_566[0:0];
  _RAND_567 = {1{`RANDOM}};
  btbV_54 = _RAND_567[0:0];
  _RAND_568 = {1{`RANDOM}};
  btbV_55 = _RAND_568[0:0];
  _RAND_569 = {1{`RANDOM}};
  btbV_56 = _RAND_569[0:0];
  _RAND_570 = {1{`RANDOM}};
  btbV_57 = _RAND_570[0:0];
  _RAND_571 = {1{`RANDOM}};
  btbV_58 = _RAND_571[0:0];
  _RAND_572 = {1{`RANDOM}};
  btbV_59 = _RAND_572[0:0];
  _RAND_573 = {1{`RANDOM}};
  btbV_60 = _RAND_573[0:0];
  _RAND_574 = {1{`RANDOM}};
  btbV_61 = _RAND_574[0:0];
  _RAND_575 = {1{`RANDOM}};
  btbV_62 = _RAND_575[0:0];
  _RAND_576 = {1{`RANDOM}};
  btbV_63 = _RAND_576[0:0];
  _RAND_577 = {1{`RANDOM}};
  btbV_64 = _RAND_577[0:0];
  _RAND_578 = {1{`RANDOM}};
  btbV_65 = _RAND_578[0:0];
  _RAND_579 = {1{`RANDOM}};
  btbV_66 = _RAND_579[0:0];
  _RAND_580 = {1{`RANDOM}};
  btbV_67 = _RAND_580[0:0];
  _RAND_581 = {1{`RANDOM}};
  btbV_68 = _RAND_581[0:0];
  _RAND_582 = {1{`RANDOM}};
  btbV_69 = _RAND_582[0:0];
  _RAND_583 = {1{`RANDOM}};
  btbV_70 = _RAND_583[0:0];
  _RAND_584 = {1{`RANDOM}};
  btbV_71 = _RAND_584[0:0];
  _RAND_585 = {1{`RANDOM}};
  btbV_72 = _RAND_585[0:0];
  _RAND_586 = {1{`RANDOM}};
  btbV_73 = _RAND_586[0:0];
  _RAND_587 = {1{`RANDOM}};
  btbV_74 = _RAND_587[0:0];
  _RAND_588 = {1{`RANDOM}};
  btbV_75 = _RAND_588[0:0];
  _RAND_589 = {1{`RANDOM}};
  btbV_76 = _RAND_589[0:0];
  _RAND_590 = {1{`RANDOM}};
  btbV_77 = _RAND_590[0:0];
  _RAND_591 = {1{`RANDOM}};
  btbV_78 = _RAND_591[0:0];
  _RAND_592 = {1{`RANDOM}};
  btbV_79 = _RAND_592[0:0];
  _RAND_593 = {1{`RANDOM}};
  btbV_80 = _RAND_593[0:0];
  _RAND_594 = {1{`RANDOM}};
  btbV_81 = _RAND_594[0:0];
  _RAND_595 = {1{`RANDOM}};
  btbV_82 = _RAND_595[0:0];
  _RAND_596 = {1{`RANDOM}};
  btbV_83 = _RAND_596[0:0];
  _RAND_597 = {1{`RANDOM}};
  btbV_84 = _RAND_597[0:0];
  _RAND_598 = {1{`RANDOM}};
  btbV_85 = _RAND_598[0:0];
  _RAND_599 = {1{`RANDOM}};
  btbV_86 = _RAND_599[0:0];
  _RAND_600 = {1{`RANDOM}};
  btbV_87 = _RAND_600[0:0];
  _RAND_601 = {1{`RANDOM}};
  btbV_88 = _RAND_601[0:0];
  _RAND_602 = {1{`RANDOM}};
  btbV_89 = _RAND_602[0:0];
  _RAND_603 = {1{`RANDOM}};
  btbV_90 = _RAND_603[0:0];
  _RAND_604 = {1{`RANDOM}};
  btbV_91 = _RAND_604[0:0];
  _RAND_605 = {1{`RANDOM}};
  btbV_92 = _RAND_605[0:0];
  _RAND_606 = {1{`RANDOM}};
  btbV_93 = _RAND_606[0:0];
  _RAND_607 = {1{`RANDOM}};
  btbV_94 = _RAND_607[0:0];
  _RAND_608 = {1{`RANDOM}};
  btbV_95 = _RAND_608[0:0];
  _RAND_609 = {1{`RANDOM}};
  btbV_96 = _RAND_609[0:0];
  _RAND_610 = {1{`RANDOM}};
  btbV_97 = _RAND_610[0:0];
  _RAND_611 = {1{`RANDOM}};
  btbV_98 = _RAND_611[0:0];
  _RAND_612 = {1{`RANDOM}};
  btbV_99 = _RAND_612[0:0];
  _RAND_613 = {1{`RANDOM}};
  btbV_100 = _RAND_613[0:0];
  _RAND_614 = {1{`RANDOM}};
  btbV_101 = _RAND_614[0:0];
  _RAND_615 = {1{`RANDOM}};
  btbV_102 = _RAND_615[0:0];
  _RAND_616 = {1{`RANDOM}};
  btbV_103 = _RAND_616[0:0];
  _RAND_617 = {1{`RANDOM}};
  btbV_104 = _RAND_617[0:0];
  _RAND_618 = {1{`RANDOM}};
  btbV_105 = _RAND_618[0:0];
  _RAND_619 = {1{`RANDOM}};
  btbV_106 = _RAND_619[0:0];
  _RAND_620 = {1{`RANDOM}};
  btbV_107 = _RAND_620[0:0];
  _RAND_621 = {1{`RANDOM}};
  btbV_108 = _RAND_621[0:0];
  _RAND_622 = {1{`RANDOM}};
  btbV_109 = _RAND_622[0:0];
  _RAND_623 = {1{`RANDOM}};
  btbV_110 = _RAND_623[0:0];
  _RAND_624 = {1{`RANDOM}};
  btbV_111 = _RAND_624[0:0];
  _RAND_625 = {1{`RANDOM}};
  btbV_112 = _RAND_625[0:0];
  _RAND_626 = {1{`RANDOM}};
  btbV_113 = _RAND_626[0:0];
  _RAND_627 = {1{`RANDOM}};
  btbV_114 = _RAND_627[0:0];
  _RAND_628 = {1{`RANDOM}};
  btbV_115 = _RAND_628[0:0];
  _RAND_629 = {1{`RANDOM}};
  btbV_116 = _RAND_629[0:0];
  _RAND_630 = {1{`RANDOM}};
  btbV_117 = _RAND_630[0:0];
  _RAND_631 = {1{`RANDOM}};
  btbV_118 = _RAND_631[0:0];
  _RAND_632 = {1{`RANDOM}};
  btbV_119 = _RAND_632[0:0];
  _RAND_633 = {1{`RANDOM}};
  btbV_120 = _RAND_633[0:0];
  _RAND_634 = {1{`RANDOM}};
  btbV_121 = _RAND_634[0:0];
  _RAND_635 = {1{`RANDOM}};
  btbV_122 = _RAND_635[0:0];
  _RAND_636 = {1{`RANDOM}};
  btbV_123 = _RAND_636[0:0];
  _RAND_637 = {1{`RANDOM}};
  btbV_124 = _RAND_637[0:0];
  _RAND_638 = {1{`RANDOM}};
  btbV_125 = _RAND_638[0:0];
  _RAND_639 = {1{`RANDOM}};
  btbV_126 = _RAND_639[0:0];
  _RAND_640 = {1{`RANDOM}};
  btbV_127 = _RAND_640[0:0];
  _RAND_641 = {1{`RANDOM}};
  btbTag_0 = _RAND_641[6:0];
  _RAND_642 = {1{`RANDOM}};
  btbTag_1 = _RAND_642[6:0];
  _RAND_643 = {1{`RANDOM}};
  btbTag_2 = _RAND_643[6:0];
  _RAND_644 = {1{`RANDOM}};
  btbTag_3 = _RAND_644[6:0];
  _RAND_645 = {1{`RANDOM}};
  btbTag_4 = _RAND_645[6:0];
  _RAND_646 = {1{`RANDOM}};
  btbTag_5 = _RAND_646[6:0];
  _RAND_647 = {1{`RANDOM}};
  btbTag_6 = _RAND_647[6:0];
  _RAND_648 = {1{`RANDOM}};
  btbTag_7 = _RAND_648[6:0];
  _RAND_649 = {1{`RANDOM}};
  btbTag_8 = _RAND_649[6:0];
  _RAND_650 = {1{`RANDOM}};
  btbTag_9 = _RAND_650[6:0];
  _RAND_651 = {1{`RANDOM}};
  btbTag_10 = _RAND_651[6:0];
  _RAND_652 = {1{`RANDOM}};
  btbTag_11 = _RAND_652[6:0];
  _RAND_653 = {1{`RANDOM}};
  btbTag_12 = _RAND_653[6:0];
  _RAND_654 = {1{`RANDOM}};
  btbTag_13 = _RAND_654[6:0];
  _RAND_655 = {1{`RANDOM}};
  btbTag_14 = _RAND_655[6:0];
  _RAND_656 = {1{`RANDOM}};
  btbTag_15 = _RAND_656[6:0];
  _RAND_657 = {1{`RANDOM}};
  btbTag_16 = _RAND_657[6:0];
  _RAND_658 = {1{`RANDOM}};
  btbTag_17 = _RAND_658[6:0];
  _RAND_659 = {1{`RANDOM}};
  btbTag_18 = _RAND_659[6:0];
  _RAND_660 = {1{`RANDOM}};
  btbTag_19 = _RAND_660[6:0];
  _RAND_661 = {1{`RANDOM}};
  btbTag_20 = _RAND_661[6:0];
  _RAND_662 = {1{`RANDOM}};
  btbTag_21 = _RAND_662[6:0];
  _RAND_663 = {1{`RANDOM}};
  btbTag_22 = _RAND_663[6:0];
  _RAND_664 = {1{`RANDOM}};
  btbTag_23 = _RAND_664[6:0];
  _RAND_665 = {1{`RANDOM}};
  btbTag_24 = _RAND_665[6:0];
  _RAND_666 = {1{`RANDOM}};
  btbTag_25 = _RAND_666[6:0];
  _RAND_667 = {1{`RANDOM}};
  btbTag_26 = _RAND_667[6:0];
  _RAND_668 = {1{`RANDOM}};
  btbTag_27 = _RAND_668[6:0];
  _RAND_669 = {1{`RANDOM}};
  btbTag_28 = _RAND_669[6:0];
  _RAND_670 = {1{`RANDOM}};
  btbTag_29 = _RAND_670[6:0];
  _RAND_671 = {1{`RANDOM}};
  btbTag_30 = _RAND_671[6:0];
  _RAND_672 = {1{`RANDOM}};
  btbTag_31 = _RAND_672[6:0];
  _RAND_673 = {1{`RANDOM}};
  btbTag_32 = _RAND_673[6:0];
  _RAND_674 = {1{`RANDOM}};
  btbTag_33 = _RAND_674[6:0];
  _RAND_675 = {1{`RANDOM}};
  btbTag_34 = _RAND_675[6:0];
  _RAND_676 = {1{`RANDOM}};
  btbTag_35 = _RAND_676[6:0];
  _RAND_677 = {1{`RANDOM}};
  btbTag_36 = _RAND_677[6:0];
  _RAND_678 = {1{`RANDOM}};
  btbTag_37 = _RAND_678[6:0];
  _RAND_679 = {1{`RANDOM}};
  btbTag_38 = _RAND_679[6:0];
  _RAND_680 = {1{`RANDOM}};
  btbTag_39 = _RAND_680[6:0];
  _RAND_681 = {1{`RANDOM}};
  btbTag_40 = _RAND_681[6:0];
  _RAND_682 = {1{`RANDOM}};
  btbTag_41 = _RAND_682[6:0];
  _RAND_683 = {1{`RANDOM}};
  btbTag_42 = _RAND_683[6:0];
  _RAND_684 = {1{`RANDOM}};
  btbTag_43 = _RAND_684[6:0];
  _RAND_685 = {1{`RANDOM}};
  btbTag_44 = _RAND_685[6:0];
  _RAND_686 = {1{`RANDOM}};
  btbTag_45 = _RAND_686[6:0];
  _RAND_687 = {1{`RANDOM}};
  btbTag_46 = _RAND_687[6:0];
  _RAND_688 = {1{`RANDOM}};
  btbTag_47 = _RAND_688[6:0];
  _RAND_689 = {1{`RANDOM}};
  btbTag_48 = _RAND_689[6:0];
  _RAND_690 = {1{`RANDOM}};
  btbTag_49 = _RAND_690[6:0];
  _RAND_691 = {1{`RANDOM}};
  btbTag_50 = _RAND_691[6:0];
  _RAND_692 = {1{`RANDOM}};
  btbTag_51 = _RAND_692[6:0];
  _RAND_693 = {1{`RANDOM}};
  btbTag_52 = _RAND_693[6:0];
  _RAND_694 = {1{`RANDOM}};
  btbTag_53 = _RAND_694[6:0];
  _RAND_695 = {1{`RANDOM}};
  btbTag_54 = _RAND_695[6:0];
  _RAND_696 = {1{`RANDOM}};
  btbTag_55 = _RAND_696[6:0];
  _RAND_697 = {1{`RANDOM}};
  btbTag_56 = _RAND_697[6:0];
  _RAND_698 = {1{`RANDOM}};
  btbTag_57 = _RAND_698[6:0];
  _RAND_699 = {1{`RANDOM}};
  btbTag_58 = _RAND_699[6:0];
  _RAND_700 = {1{`RANDOM}};
  btbTag_59 = _RAND_700[6:0];
  _RAND_701 = {1{`RANDOM}};
  btbTag_60 = _RAND_701[6:0];
  _RAND_702 = {1{`RANDOM}};
  btbTag_61 = _RAND_702[6:0];
  _RAND_703 = {1{`RANDOM}};
  btbTag_62 = _RAND_703[6:0];
  _RAND_704 = {1{`RANDOM}};
  btbTag_63 = _RAND_704[6:0];
  _RAND_705 = {1{`RANDOM}};
  btbTag_64 = _RAND_705[6:0];
  _RAND_706 = {1{`RANDOM}};
  btbTag_65 = _RAND_706[6:0];
  _RAND_707 = {1{`RANDOM}};
  btbTag_66 = _RAND_707[6:0];
  _RAND_708 = {1{`RANDOM}};
  btbTag_67 = _RAND_708[6:0];
  _RAND_709 = {1{`RANDOM}};
  btbTag_68 = _RAND_709[6:0];
  _RAND_710 = {1{`RANDOM}};
  btbTag_69 = _RAND_710[6:0];
  _RAND_711 = {1{`RANDOM}};
  btbTag_70 = _RAND_711[6:0];
  _RAND_712 = {1{`RANDOM}};
  btbTag_71 = _RAND_712[6:0];
  _RAND_713 = {1{`RANDOM}};
  btbTag_72 = _RAND_713[6:0];
  _RAND_714 = {1{`RANDOM}};
  btbTag_73 = _RAND_714[6:0];
  _RAND_715 = {1{`RANDOM}};
  btbTag_74 = _RAND_715[6:0];
  _RAND_716 = {1{`RANDOM}};
  btbTag_75 = _RAND_716[6:0];
  _RAND_717 = {1{`RANDOM}};
  btbTag_76 = _RAND_717[6:0];
  _RAND_718 = {1{`RANDOM}};
  btbTag_77 = _RAND_718[6:0];
  _RAND_719 = {1{`RANDOM}};
  btbTag_78 = _RAND_719[6:0];
  _RAND_720 = {1{`RANDOM}};
  btbTag_79 = _RAND_720[6:0];
  _RAND_721 = {1{`RANDOM}};
  btbTag_80 = _RAND_721[6:0];
  _RAND_722 = {1{`RANDOM}};
  btbTag_81 = _RAND_722[6:0];
  _RAND_723 = {1{`RANDOM}};
  btbTag_82 = _RAND_723[6:0];
  _RAND_724 = {1{`RANDOM}};
  btbTag_83 = _RAND_724[6:0];
  _RAND_725 = {1{`RANDOM}};
  btbTag_84 = _RAND_725[6:0];
  _RAND_726 = {1{`RANDOM}};
  btbTag_85 = _RAND_726[6:0];
  _RAND_727 = {1{`RANDOM}};
  btbTag_86 = _RAND_727[6:0];
  _RAND_728 = {1{`RANDOM}};
  btbTag_87 = _RAND_728[6:0];
  _RAND_729 = {1{`RANDOM}};
  btbTag_88 = _RAND_729[6:0];
  _RAND_730 = {1{`RANDOM}};
  btbTag_89 = _RAND_730[6:0];
  _RAND_731 = {1{`RANDOM}};
  btbTag_90 = _RAND_731[6:0];
  _RAND_732 = {1{`RANDOM}};
  btbTag_91 = _RAND_732[6:0];
  _RAND_733 = {1{`RANDOM}};
  btbTag_92 = _RAND_733[6:0];
  _RAND_734 = {1{`RANDOM}};
  btbTag_93 = _RAND_734[6:0];
  _RAND_735 = {1{`RANDOM}};
  btbTag_94 = _RAND_735[6:0];
  _RAND_736 = {1{`RANDOM}};
  btbTag_95 = _RAND_736[6:0];
  _RAND_737 = {1{`RANDOM}};
  btbTag_96 = _RAND_737[6:0];
  _RAND_738 = {1{`RANDOM}};
  btbTag_97 = _RAND_738[6:0];
  _RAND_739 = {1{`RANDOM}};
  btbTag_98 = _RAND_739[6:0];
  _RAND_740 = {1{`RANDOM}};
  btbTag_99 = _RAND_740[6:0];
  _RAND_741 = {1{`RANDOM}};
  btbTag_100 = _RAND_741[6:0];
  _RAND_742 = {1{`RANDOM}};
  btbTag_101 = _RAND_742[6:0];
  _RAND_743 = {1{`RANDOM}};
  btbTag_102 = _RAND_743[6:0];
  _RAND_744 = {1{`RANDOM}};
  btbTag_103 = _RAND_744[6:0];
  _RAND_745 = {1{`RANDOM}};
  btbTag_104 = _RAND_745[6:0];
  _RAND_746 = {1{`RANDOM}};
  btbTag_105 = _RAND_746[6:0];
  _RAND_747 = {1{`RANDOM}};
  btbTag_106 = _RAND_747[6:0];
  _RAND_748 = {1{`RANDOM}};
  btbTag_107 = _RAND_748[6:0];
  _RAND_749 = {1{`RANDOM}};
  btbTag_108 = _RAND_749[6:0];
  _RAND_750 = {1{`RANDOM}};
  btbTag_109 = _RAND_750[6:0];
  _RAND_751 = {1{`RANDOM}};
  btbTag_110 = _RAND_751[6:0];
  _RAND_752 = {1{`RANDOM}};
  btbTag_111 = _RAND_752[6:0];
  _RAND_753 = {1{`RANDOM}};
  btbTag_112 = _RAND_753[6:0];
  _RAND_754 = {1{`RANDOM}};
  btbTag_113 = _RAND_754[6:0];
  _RAND_755 = {1{`RANDOM}};
  btbTag_114 = _RAND_755[6:0];
  _RAND_756 = {1{`RANDOM}};
  btbTag_115 = _RAND_756[6:0];
  _RAND_757 = {1{`RANDOM}};
  btbTag_116 = _RAND_757[6:0];
  _RAND_758 = {1{`RANDOM}};
  btbTag_117 = _RAND_758[6:0];
  _RAND_759 = {1{`RANDOM}};
  btbTag_118 = _RAND_759[6:0];
  _RAND_760 = {1{`RANDOM}};
  btbTag_119 = _RAND_760[6:0];
  _RAND_761 = {1{`RANDOM}};
  btbTag_120 = _RAND_761[6:0];
  _RAND_762 = {1{`RANDOM}};
  btbTag_121 = _RAND_762[6:0];
  _RAND_763 = {1{`RANDOM}};
  btbTag_122 = _RAND_763[6:0];
  _RAND_764 = {1{`RANDOM}};
  btbTag_123 = _RAND_764[6:0];
  _RAND_765 = {1{`RANDOM}};
  btbTag_124 = _RAND_765[6:0];
  _RAND_766 = {1{`RANDOM}};
  btbTag_125 = _RAND_766[6:0];
  _RAND_767 = {1{`RANDOM}};
  btbTag_126 = _RAND_767[6:0];
  _RAND_768 = {1{`RANDOM}};
  btbTag_127 = _RAND_768[6:0];
  _RAND_769 = {1{`RANDOM}};
  btbMeta_0 = _RAND_769[31:0];
  _RAND_770 = {1{`RANDOM}};
  btbMeta_1 = _RAND_770[31:0];
  _RAND_771 = {1{`RANDOM}};
  btbMeta_2 = _RAND_771[31:0];
  _RAND_772 = {1{`RANDOM}};
  btbMeta_3 = _RAND_772[31:0];
  _RAND_773 = {1{`RANDOM}};
  btbMeta_4 = _RAND_773[31:0];
  _RAND_774 = {1{`RANDOM}};
  btbMeta_5 = _RAND_774[31:0];
  _RAND_775 = {1{`RANDOM}};
  btbMeta_6 = _RAND_775[31:0];
  _RAND_776 = {1{`RANDOM}};
  btbMeta_7 = _RAND_776[31:0];
  _RAND_777 = {1{`RANDOM}};
  btbMeta_8 = _RAND_777[31:0];
  _RAND_778 = {1{`RANDOM}};
  btbMeta_9 = _RAND_778[31:0];
  _RAND_779 = {1{`RANDOM}};
  btbMeta_10 = _RAND_779[31:0];
  _RAND_780 = {1{`RANDOM}};
  btbMeta_11 = _RAND_780[31:0];
  _RAND_781 = {1{`RANDOM}};
  btbMeta_12 = _RAND_781[31:0];
  _RAND_782 = {1{`RANDOM}};
  btbMeta_13 = _RAND_782[31:0];
  _RAND_783 = {1{`RANDOM}};
  btbMeta_14 = _RAND_783[31:0];
  _RAND_784 = {1{`RANDOM}};
  btbMeta_15 = _RAND_784[31:0];
  _RAND_785 = {1{`RANDOM}};
  btbMeta_16 = _RAND_785[31:0];
  _RAND_786 = {1{`RANDOM}};
  btbMeta_17 = _RAND_786[31:0];
  _RAND_787 = {1{`RANDOM}};
  btbMeta_18 = _RAND_787[31:0];
  _RAND_788 = {1{`RANDOM}};
  btbMeta_19 = _RAND_788[31:0];
  _RAND_789 = {1{`RANDOM}};
  btbMeta_20 = _RAND_789[31:0];
  _RAND_790 = {1{`RANDOM}};
  btbMeta_21 = _RAND_790[31:0];
  _RAND_791 = {1{`RANDOM}};
  btbMeta_22 = _RAND_791[31:0];
  _RAND_792 = {1{`RANDOM}};
  btbMeta_23 = _RAND_792[31:0];
  _RAND_793 = {1{`RANDOM}};
  btbMeta_24 = _RAND_793[31:0];
  _RAND_794 = {1{`RANDOM}};
  btbMeta_25 = _RAND_794[31:0];
  _RAND_795 = {1{`RANDOM}};
  btbMeta_26 = _RAND_795[31:0];
  _RAND_796 = {1{`RANDOM}};
  btbMeta_27 = _RAND_796[31:0];
  _RAND_797 = {1{`RANDOM}};
  btbMeta_28 = _RAND_797[31:0];
  _RAND_798 = {1{`RANDOM}};
  btbMeta_29 = _RAND_798[31:0];
  _RAND_799 = {1{`RANDOM}};
  btbMeta_30 = _RAND_799[31:0];
  _RAND_800 = {1{`RANDOM}};
  btbMeta_31 = _RAND_800[31:0];
  _RAND_801 = {1{`RANDOM}};
  btbMeta_32 = _RAND_801[31:0];
  _RAND_802 = {1{`RANDOM}};
  btbMeta_33 = _RAND_802[31:0];
  _RAND_803 = {1{`RANDOM}};
  btbMeta_34 = _RAND_803[31:0];
  _RAND_804 = {1{`RANDOM}};
  btbMeta_35 = _RAND_804[31:0];
  _RAND_805 = {1{`RANDOM}};
  btbMeta_36 = _RAND_805[31:0];
  _RAND_806 = {1{`RANDOM}};
  btbMeta_37 = _RAND_806[31:0];
  _RAND_807 = {1{`RANDOM}};
  btbMeta_38 = _RAND_807[31:0];
  _RAND_808 = {1{`RANDOM}};
  btbMeta_39 = _RAND_808[31:0];
  _RAND_809 = {1{`RANDOM}};
  btbMeta_40 = _RAND_809[31:0];
  _RAND_810 = {1{`RANDOM}};
  btbMeta_41 = _RAND_810[31:0];
  _RAND_811 = {1{`RANDOM}};
  btbMeta_42 = _RAND_811[31:0];
  _RAND_812 = {1{`RANDOM}};
  btbMeta_43 = _RAND_812[31:0];
  _RAND_813 = {1{`RANDOM}};
  btbMeta_44 = _RAND_813[31:0];
  _RAND_814 = {1{`RANDOM}};
  btbMeta_45 = _RAND_814[31:0];
  _RAND_815 = {1{`RANDOM}};
  btbMeta_46 = _RAND_815[31:0];
  _RAND_816 = {1{`RANDOM}};
  btbMeta_47 = _RAND_816[31:0];
  _RAND_817 = {1{`RANDOM}};
  btbMeta_48 = _RAND_817[31:0];
  _RAND_818 = {1{`RANDOM}};
  btbMeta_49 = _RAND_818[31:0];
  _RAND_819 = {1{`RANDOM}};
  btbMeta_50 = _RAND_819[31:0];
  _RAND_820 = {1{`RANDOM}};
  btbMeta_51 = _RAND_820[31:0];
  _RAND_821 = {1{`RANDOM}};
  btbMeta_52 = _RAND_821[31:0];
  _RAND_822 = {1{`RANDOM}};
  btbMeta_53 = _RAND_822[31:0];
  _RAND_823 = {1{`RANDOM}};
  btbMeta_54 = _RAND_823[31:0];
  _RAND_824 = {1{`RANDOM}};
  btbMeta_55 = _RAND_824[31:0];
  _RAND_825 = {1{`RANDOM}};
  btbMeta_56 = _RAND_825[31:0];
  _RAND_826 = {1{`RANDOM}};
  btbMeta_57 = _RAND_826[31:0];
  _RAND_827 = {1{`RANDOM}};
  btbMeta_58 = _RAND_827[31:0];
  _RAND_828 = {1{`RANDOM}};
  btbMeta_59 = _RAND_828[31:0];
  _RAND_829 = {1{`RANDOM}};
  btbMeta_60 = _RAND_829[31:0];
  _RAND_830 = {1{`RANDOM}};
  btbMeta_61 = _RAND_830[31:0];
  _RAND_831 = {1{`RANDOM}};
  btbMeta_62 = _RAND_831[31:0];
  _RAND_832 = {1{`RANDOM}};
  btbMeta_63 = _RAND_832[31:0];
  _RAND_833 = {1{`RANDOM}};
  btbMeta_64 = _RAND_833[31:0];
  _RAND_834 = {1{`RANDOM}};
  btbMeta_65 = _RAND_834[31:0];
  _RAND_835 = {1{`RANDOM}};
  btbMeta_66 = _RAND_835[31:0];
  _RAND_836 = {1{`RANDOM}};
  btbMeta_67 = _RAND_836[31:0];
  _RAND_837 = {1{`RANDOM}};
  btbMeta_68 = _RAND_837[31:0];
  _RAND_838 = {1{`RANDOM}};
  btbMeta_69 = _RAND_838[31:0];
  _RAND_839 = {1{`RANDOM}};
  btbMeta_70 = _RAND_839[31:0];
  _RAND_840 = {1{`RANDOM}};
  btbMeta_71 = _RAND_840[31:0];
  _RAND_841 = {1{`RANDOM}};
  btbMeta_72 = _RAND_841[31:0];
  _RAND_842 = {1{`RANDOM}};
  btbMeta_73 = _RAND_842[31:0];
  _RAND_843 = {1{`RANDOM}};
  btbMeta_74 = _RAND_843[31:0];
  _RAND_844 = {1{`RANDOM}};
  btbMeta_75 = _RAND_844[31:0];
  _RAND_845 = {1{`RANDOM}};
  btbMeta_76 = _RAND_845[31:0];
  _RAND_846 = {1{`RANDOM}};
  btbMeta_77 = _RAND_846[31:0];
  _RAND_847 = {1{`RANDOM}};
  btbMeta_78 = _RAND_847[31:0];
  _RAND_848 = {1{`RANDOM}};
  btbMeta_79 = _RAND_848[31:0];
  _RAND_849 = {1{`RANDOM}};
  btbMeta_80 = _RAND_849[31:0];
  _RAND_850 = {1{`RANDOM}};
  btbMeta_81 = _RAND_850[31:0];
  _RAND_851 = {1{`RANDOM}};
  btbMeta_82 = _RAND_851[31:0];
  _RAND_852 = {1{`RANDOM}};
  btbMeta_83 = _RAND_852[31:0];
  _RAND_853 = {1{`RANDOM}};
  btbMeta_84 = _RAND_853[31:0];
  _RAND_854 = {1{`RANDOM}};
  btbMeta_85 = _RAND_854[31:0];
  _RAND_855 = {1{`RANDOM}};
  btbMeta_86 = _RAND_855[31:0];
  _RAND_856 = {1{`RANDOM}};
  btbMeta_87 = _RAND_856[31:0];
  _RAND_857 = {1{`RANDOM}};
  btbMeta_88 = _RAND_857[31:0];
  _RAND_858 = {1{`RANDOM}};
  btbMeta_89 = _RAND_858[31:0];
  _RAND_859 = {1{`RANDOM}};
  btbMeta_90 = _RAND_859[31:0];
  _RAND_860 = {1{`RANDOM}};
  btbMeta_91 = _RAND_860[31:0];
  _RAND_861 = {1{`RANDOM}};
  btbMeta_92 = _RAND_861[31:0];
  _RAND_862 = {1{`RANDOM}};
  btbMeta_93 = _RAND_862[31:0];
  _RAND_863 = {1{`RANDOM}};
  btbMeta_94 = _RAND_863[31:0];
  _RAND_864 = {1{`RANDOM}};
  btbMeta_95 = _RAND_864[31:0];
  _RAND_865 = {1{`RANDOM}};
  btbMeta_96 = _RAND_865[31:0];
  _RAND_866 = {1{`RANDOM}};
  btbMeta_97 = _RAND_866[31:0];
  _RAND_867 = {1{`RANDOM}};
  btbMeta_98 = _RAND_867[31:0];
  _RAND_868 = {1{`RANDOM}};
  btbMeta_99 = _RAND_868[31:0];
  _RAND_869 = {1{`RANDOM}};
  btbMeta_100 = _RAND_869[31:0];
  _RAND_870 = {1{`RANDOM}};
  btbMeta_101 = _RAND_870[31:0];
  _RAND_871 = {1{`RANDOM}};
  btbMeta_102 = _RAND_871[31:0];
  _RAND_872 = {1{`RANDOM}};
  btbMeta_103 = _RAND_872[31:0];
  _RAND_873 = {1{`RANDOM}};
  btbMeta_104 = _RAND_873[31:0];
  _RAND_874 = {1{`RANDOM}};
  btbMeta_105 = _RAND_874[31:0];
  _RAND_875 = {1{`RANDOM}};
  btbMeta_106 = _RAND_875[31:0];
  _RAND_876 = {1{`RANDOM}};
  btbMeta_107 = _RAND_876[31:0];
  _RAND_877 = {1{`RANDOM}};
  btbMeta_108 = _RAND_877[31:0];
  _RAND_878 = {1{`RANDOM}};
  btbMeta_109 = _RAND_878[31:0];
  _RAND_879 = {1{`RANDOM}};
  btbMeta_110 = _RAND_879[31:0];
  _RAND_880 = {1{`RANDOM}};
  btbMeta_111 = _RAND_880[31:0];
  _RAND_881 = {1{`RANDOM}};
  btbMeta_112 = _RAND_881[31:0];
  _RAND_882 = {1{`RANDOM}};
  btbMeta_113 = _RAND_882[31:0];
  _RAND_883 = {1{`RANDOM}};
  btbMeta_114 = _RAND_883[31:0];
  _RAND_884 = {1{`RANDOM}};
  btbMeta_115 = _RAND_884[31:0];
  _RAND_885 = {1{`RANDOM}};
  btbMeta_116 = _RAND_885[31:0];
  _RAND_886 = {1{`RANDOM}};
  btbMeta_117 = _RAND_886[31:0];
  _RAND_887 = {1{`RANDOM}};
  btbMeta_118 = _RAND_887[31:0];
  _RAND_888 = {1{`RANDOM}};
  btbMeta_119 = _RAND_888[31:0];
  _RAND_889 = {1{`RANDOM}};
  btbMeta_120 = _RAND_889[31:0];
  _RAND_890 = {1{`RANDOM}};
  btbMeta_121 = _RAND_890[31:0];
  _RAND_891 = {1{`RANDOM}};
  btbMeta_122 = _RAND_891[31:0];
  _RAND_892 = {1{`RANDOM}};
  btbMeta_123 = _RAND_892[31:0];
  _RAND_893 = {1{`RANDOM}};
  btbMeta_124 = _RAND_893[31:0];
  _RAND_894 = {1{`RANDOM}};
  btbMeta_125 = _RAND_894[31:0];
  _RAND_895 = {1{`RANDOM}};
  btbMeta_126 = _RAND_895[31:0];
  _RAND_896 = {1{`RANDOM}};
  btbMeta_127 = _RAND_896[31:0];
  _RAND_897 = {1{`RANDOM}};
  io_ready_REG = _RAND_897[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module InstFetch(
  input         clock,
  input         reset,
  output        io_imem_inst_valid,
  input         io_imem_inst_ready,
  output [31:0] io_imem_inst_addr,
  input  [31:0] io_imem_inst_read,
  input         io_takenValid,
  input         io_takenValidJalr,
  input         io_takenMiss,
  input         io_exTakenPre,
  input  [31:0] io_takenPC,
  input  [31:0] io_nextPC,
  input         io_stall,
  input         io_exc,
  input         io_intr,
  output        io_out_valid,
  output [31:0] io_out_pc,
  output [31:0] io_out_inst,
  output        io_out_takenPre,
  output [31:0] io_out_takenPrePC,
  output        io_IFDone,
  output        io_preRs1En,
  output [4:0]  io_preRs1Addr,
  input  [63:0] io_preRs1Data,
  input  [63:0] io_preRs1x1Data,
  input         io_exeX1En,
  input  [63:0] io_exeAluRes,
  input         io_memX1En,
  input  [63:0] io_memAluRes,
  input         io_wbRdEn,
  input  [4:0]  io_wbRdAddr,
  input  [63:0] io_wbRdData
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] minidec_io_inst; // @[InstFetch.scala 50:23]
  wire  minidec_io_rs1En; // @[InstFetch.scala 50:23]
  wire [4:0] minidec_io_rs1Addr; // @[InstFetch.scala 50:23]
  wire  minidec_io_bjp; // @[InstFetch.scala 50:23]
  wire  minidec_io_jal; // @[InstFetch.scala 50:23]
  wire  minidec_io_jalr; // @[InstFetch.scala 50:23]
  wire  minidec_io_bxx; // @[InstFetch.scala 50:23]
  wire [63:0] minidec_io_imm; // @[InstFetch.scala 50:23]
  wire  bht_clock; // @[InstFetch.scala 51:19]
  wire  bht_reset; // @[InstFetch.scala 51:19]
  wire  bht_io_valid; // @[InstFetch.scala 51:19]
  wire  bht_io_fire; // @[InstFetch.scala 51:19]
  wire [31:0] bht_io_pc; // @[InstFetch.scala 51:19]
  wire  bht_io_jal; // @[InstFetch.scala 51:19]
  wire  bht_io_jalr; // @[InstFetch.scala 51:19]
  wire  bht_io_bxx; // @[InstFetch.scala 51:19]
  wire [63:0] bht_io_imm; // @[InstFetch.scala 51:19]
  wire [4:0] bht_io_rs1Addr; // @[InstFetch.scala 51:19]
  wire [63:0] bht_io_rs1Data; // @[InstFetch.scala 51:19]
  wire [63:0] bht_io_rs1x1Data; // @[InstFetch.scala 51:19]
  wire  bht_io_exeX1En; // @[InstFetch.scala 51:19]
  wire [63:0] bht_io_exeAluRes; // @[InstFetch.scala 51:19]
  wire  bht_io_memX1En; // @[InstFetch.scala 51:19]
  wire [63:0] bht_io_memAluRes; // @[InstFetch.scala 51:19]
  wire  bht_io_wbRdEn; // @[InstFetch.scala 51:19]
  wire [4:0] bht_io_wbRdAddr; // @[InstFetch.scala 51:19]
  wire [63:0] bht_io_wbRdData; // @[InstFetch.scala 51:19]
  wire  bht_io_takenValid; // @[InstFetch.scala 51:19]
  wire  bht_io_takenValidJalr; // @[InstFetch.scala 51:19]
  wire  bht_io_takenMiss; // @[InstFetch.scala 51:19]
  wire  bht_io_exTakenPre; // @[InstFetch.scala 51:19]
  wire [31:0] bht_io_takenPC; // @[InstFetch.scala 51:19]
  wire [31:0] bht_io_nextPC; // @[InstFetch.scala 51:19]
  wire  bht_io_takenPre; // @[InstFetch.scala 51:19]
  wire [31:0] bht_io_takenPrePC; // @[InstFetch.scala 51:19]
  wire  bht_io_ready; // @[InstFetch.scala 51:19]
  reg [31:0] pc; // @[InstFetch.scala 53:19]
  reg [31:0] inst; // @[InstFetch.scala 54:21]
  wire  _io_imem_inst_valid_T = ~io_stall; // @[InstFetch.scala 57:25]
  wire  fire = io_imem_inst_valid & io_imem_inst_ready; // @[InstFetch.scala 62:33]
  wire  ifPcEn = bht_io_ready & _io_imem_inst_valid_T & ~io_intr; // @[InstFetch.scala 67:37]
  wire [31:0] _ifPC_T_3 = pc + 32'h4; // @[InstFetch.scala 70:79]
  minidec minidec ( // @[InstFetch.scala 50:23]
    .io_inst(minidec_io_inst),
    .io_rs1En(minidec_io_rs1En),
    .io_rs1Addr(minidec_io_rs1Addr),
    .io_bjp(minidec_io_bjp),
    .io_jal(minidec_io_jal),
    .io_jalr(minidec_io_jalr),
    .io_bxx(minidec_io_bxx),
    .io_imm(minidec_io_imm)
  );
  bht bht ( // @[InstFetch.scala 51:19]
    .clock(bht_clock),
    .reset(bht_reset),
    .io_valid(bht_io_valid),
    .io_fire(bht_io_fire),
    .io_pc(bht_io_pc),
    .io_jal(bht_io_jal),
    .io_jalr(bht_io_jalr),
    .io_bxx(bht_io_bxx),
    .io_imm(bht_io_imm),
    .io_rs1Addr(bht_io_rs1Addr),
    .io_rs1Data(bht_io_rs1Data),
    .io_rs1x1Data(bht_io_rs1x1Data),
    .io_exeX1En(bht_io_exeX1En),
    .io_exeAluRes(bht_io_exeAluRes),
    .io_memX1En(bht_io_memX1En),
    .io_memAluRes(bht_io_memAluRes),
    .io_wbRdEn(bht_io_wbRdEn),
    .io_wbRdAddr(bht_io_wbRdAddr),
    .io_wbRdData(bht_io_wbRdData),
    .io_takenValid(bht_io_takenValid),
    .io_takenValidJalr(bht_io_takenValidJalr),
    .io_takenMiss(bht_io_takenMiss),
    .io_exTakenPre(bht_io_exTakenPre),
    .io_takenPC(bht_io_takenPC),
    .io_nextPC(bht_io_nextPC),
    .io_takenPre(bht_io_takenPre),
    .io_takenPrePC(bht_io_takenPrePC),
    .io_ready(bht_io_ready)
  );
  assign io_imem_inst_valid = ~io_stall; // @[InstFetch.scala 57:25]
  assign io_imem_inst_addr = pc; // @[InstFetch.scala 59:21]
  assign io_out_valid = bht_io_ready; // @[InstFetch.scala 110:19]
  assign io_out_pc = pc; // @[InstFetch.scala 111:19]
  assign io_out_inst = minidec_io_bxx ? inst : io_imem_inst_read; // @[InstFetch.scala 108:19]
  assign io_out_takenPre = bht_io_takenPre; // @[InstFetch.scala 133:19]
  assign io_out_takenPrePC = bht_io_takenPrePC; // @[InstFetch.scala 134:21]
  assign io_IFDone = io_stall | bht_io_ready; // @[InstFetch.scala 76:19]
  assign io_preRs1En = minidec_io_rs1En; // @[InstFetch.scala 105:15]
  assign io_preRs1Addr = minidec_io_rs1Addr; // @[InstFetch.scala 106:17]
  assign minidec_io_inst = fire & _io_imem_inst_valid_T ? io_imem_inst_read : inst; // @[InstFetch.scala 66:19]
  assign bht_clock = clock;
  assign bht_reset = reset;
  assign bht_io_valid = minidec_io_bjp; // @[InstFetch.scala 81:16]
  assign bht_io_fire = io_imem_inst_valid & io_imem_inst_ready; // @[InstFetch.scala 62:33]
  assign bht_io_pc = pc; // @[InstFetch.scala 80:13]
  assign bht_io_jal = minidec_io_jal; // @[InstFetch.scala 83:14]
  assign bht_io_jalr = minidec_io_jalr; // @[InstFetch.scala 84:15]
  assign bht_io_bxx = minidec_io_bxx; // @[InstFetch.scala 85:14]
  assign bht_io_imm = minidec_io_imm; // @[InstFetch.scala 86:14]
  assign bht_io_rs1Addr = minidec_io_rs1Addr; // @[InstFetch.scala 87:18]
  assign bht_io_rs1Data = io_preRs1Data; // @[InstFetch.scala 95:18]
  assign bht_io_rs1x1Data = io_preRs1x1Data; // @[InstFetch.scala 96:20]
  assign bht_io_exeX1En = io_exeX1En; // @[InstFetch.scala 97:18]
  assign bht_io_exeAluRes = io_exeAluRes; // @[InstFetch.scala 98:20]
  assign bht_io_memX1En = io_memX1En; // @[InstFetch.scala 99:18]
  assign bht_io_memAluRes = io_memAluRes; // @[InstFetch.scala 100:20]
  assign bht_io_wbRdEn = io_wbRdEn; // @[InstFetch.scala 101:17]
  assign bht_io_wbRdAddr = io_wbRdAddr; // @[InstFetch.scala 102:19]
  assign bht_io_wbRdData = io_wbRdData; // @[InstFetch.scala 103:19]
  assign bht_io_takenValid = io_takenValid; // @[InstFetch.scala 89:21]
  assign bht_io_takenValidJalr = io_takenValidJalr; // @[InstFetch.scala 90:25]
  assign bht_io_takenMiss = io_takenMiss; // @[InstFetch.scala 91:20]
  assign bht_io_exTakenPre = io_exTakenPre; // @[InstFetch.scala 92:21]
  assign bht_io_takenPC = io_takenPC; // @[InstFetch.scala 93:18]
  assign bht_io_nextPC = io_nextPC; // @[InstFetch.scala 94:17]
  always @(posedge clock) begin
    if (reset) begin // @[InstFetch.scala 53:19]
      pc <= 32'h80000000; // @[InstFetch.scala 53:19]
    end else if (ifPcEn) begin // @[InstFetch.scala 68:17]
      if (io_exc | io_takenMiss) begin // @[InstFetch.scala 69:20]
        pc <= io_nextPC;
      end else if (bht_io_takenPre & minidec_io_bjp) begin // @[InstFetch.scala 70:22]
        pc <= bht_io_takenPrePC;
      end else begin
        pc <= _ifPC_T_3;
      end
    end else if (io_intr) begin // @[InstFetch.scala 71:20]
      pc <= io_nextPC;
    end
    if (reset) begin // @[InstFetch.scala 54:21]
      inst <= 32'h0; // @[InstFetch.scala 54:21]
    end else if (fire & _io_imem_inst_valid_T) begin // @[InstFetch.scala 66:19]
      inst <= io_imem_inst_read;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  pc = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  inst = _RAND_1[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PipelineReg(
  input         clock,
  input         reset,
  input         io_in_valid,
  input  [31:0] io_in_pc,
  input  [31:0] io_in_inst,
  input         io_in_typeL,
  input         io_in_aluA,
  input  [1:0]  io_in_aluB,
  input  [3:0]  io_in_aluOp,
  input  [2:0]  io_in_branch,
  input  [1:0]  io_in_memtoReg,
  input         io_in_memWr,
  input  [2:0]  io_in_memOp,
  input  [31:0] io_in_memAddr,
  input         io_in_rdEn,
  input  [4:0]  io_in_rdAddr,
  input  [63:0] io_in_rs1Data,
  input  [63:0] io_in_rs2Data,
  input  [63:0] io_in_imm,
  input  [63:0] io_in_aluRes,
  input  [63:0] io_in_memData,
  input  [3:0]  io_in_csrOp,
  input         io_in_takenPre,
  input  [31:0] io_in_takenPrePC,
  output        io_out_valid,
  output [31:0] io_out_pc,
  output [31:0] io_out_inst,
  output        io_out_typeL,
  output        io_out_aluA,
  output [1:0]  io_out_aluB,
  output [3:0]  io_out_aluOp,
  output [2:0]  io_out_branch,
  output [1:0]  io_out_memtoReg,
  output        io_out_memWr,
  output [2:0]  io_out_memOp,
  output [31:0] io_out_memAddr,
  output        io_out_rdEn,
  output [4:0]  io_out_rdAddr,
  output [63:0] io_out_rs1Data,
  output [63:0] io_out_rs2Data,
  output [63:0] io_out_imm,
  output [63:0] io_out_aluRes,
  output [63:0] io_out_memData,
  output [3:0]  io_out_csrOp,
  output        io_out_takenPre,
  output [31:0] io_out_takenPrePC,
  input         io_flush,
  input         io_stall
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
`endif // RANDOMIZE_REG_INIT
  reg  reg_valid; // @[PipelineReg.scala 82:20]
  reg [31:0] reg_pc; // @[PipelineReg.scala 82:20]
  reg [31:0] reg_inst; // @[PipelineReg.scala 82:20]
  reg  reg_typeL; // @[PipelineReg.scala 82:20]
  reg  reg_aluA; // @[PipelineReg.scala 82:20]
  reg [1:0] reg_aluB; // @[PipelineReg.scala 82:20]
  reg [3:0] reg_aluOp; // @[PipelineReg.scala 82:20]
  reg [2:0] reg_branch; // @[PipelineReg.scala 82:20]
  reg [1:0] reg_memtoReg; // @[PipelineReg.scala 82:20]
  reg  reg_memWr; // @[PipelineReg.scala 82:20]
  reg [2:0] reg_memOp; // @[PipelineReg.scala 82:20]
  reg [31:0] reg_memAddr; // @[PipelineReg.scala 82:20]
  reg  reg_rdEn; // @[PipelineReg.scala 82:20]
  reg [4:0] reg_rdAddr; // @[PipelineReg.scala 82:20]
  reg [63:0] reg_rs1Data; // @[PipelineReg.scala 82:20]
  reg [63:0] reg_rs2Data; // @[PipelineReg.scala 82:20]
  reg [63:0] reg_imm; // @[PipelineReg.scala 82:20]
  reg [63:0] reg_aluRes; // @[PipelineReg.scala 82:20]
  reg [63:0] reg_memData; // @[PipelineReg.scala 82:20]
  reg [3:0] reg_csrOp; // @[PipelineReg.scala 82:20]
  reg  reg_takenPre; // @[PipelineReg.scala 82:20]
  reg [31:0] reg_takenPrePC; // @[PipelineReg.scala 82:20]
  wire  _T = ~io_stall; // @[PipelineReg.scala 84:33]
  assign io_out_valid = reg_valid; // @[PipelineReg.scala 90:10]
  assign io_out_pc = reg_pc; // @[PipelineReg.scala 90:10]
  assign io_out_inst = reg_inst; // @[PipelineReg.scala 90:10]
  assign io_out_typeL = reg_typeL; // @[PipelineReg.scala 90:10]
  assign io_out_aluA = reg_aluA; // @[PipelineReg.scala 90:10]
  assign io_out_aluB = reg_aluB; // @[PipelineReg.scala 90:10]
  assign io_out_aluOp = reg_aluOp; // @[PipelineReg.scala 90:10]
  assign io_out_branch = reg_branch; // @[PipelineReg.scala 90:10]
  assign io_out_memtoReg = reg_memtoReg; // @[PipelineReg.scala 90:10]
  assign io_out_memWr = reg_memWr; // @[PipelineReg.scala 90:10]
  assign io_out_memOp = reg_memOp; // @[PipelineReg.scala 90:10]
  assign io_out_memAddr = reg_memAddr; // @[PipelineReg.scala 90:10]
  assign io_out_rdEn = reg_rdEn; // @[PipelineReg.scala 90:10]
  assign io_out_rdAddr = reg_rdAddr; // @[PipelineReg.scala 90:10]
  assign io_out_rs1Data = reg_rs1Data; // @[PipelineReg.scala 90:10]
  assign io_out_rs2Data = reg_rs2Data; // @[PipelineReg.scala 90:10]
  assign io_out_imm = reg_imm; // @[PipelineReg.scala 90:10]
  assign io_out_aluRes = reg_aluRes; // @[PipelineReg.scala 90:10]
  assign io_out_memData = reg_memData; // @[PipelineReg.scala 90:10]
  assign io_out_csrOp = reg_csrOp; // @[PipelineReg.scala 90:10]
  assign io_out_takenPre = reg_takenPre; // @[PipelineReg.scala 90:10]
  assign io_out_takenPrePC = reg_takenPrePC; // @[PipelineReg.scala 90:10]
  always @(posedge clock) begin
    if (reset) begin // @[PipelineReg.scala 82:20]
      reg_valid <= 1'h0; // @[PipelineReg.scala 82:20]
    end else if (io_flush & ~io_stall) begin // @[PipelineReg.scala 84:44]
      reg_valid <= 1'h0; // @[PipelineReg.scala 37:14]
    end else if (_T) begin // @[PipelineReg.scala 86:27]
      reg_valid <= io_in_valid; // @[PipelineReg.scala 87:9]
    end
    if (reset) begin // @[PipelineReg.scala 82:20]
      reg_pc <= 32'h0; // @[PipelineReg.scala 82:20]
    end else if (io_flush & ~io_stall) begin // @[PipelineReg.scala 84:44]
      reg_pc <= 32'h0; // @[PipelineReg.scala 38:14]
    end else if (_T) begin // @[PipelineReg.scala 86:27]
      reg_pc <= io_in_pc; // @[PipelineReg.scala 87:9]
    end
    if (reset) begin // @[PipelineReg.scala 82:20]
      reg_inst <= 32'h0; // @[PipelineReg.scala 82:20]
    end else if (io_flush & ~io_stall) begin // @[PipelineReg.scala 84:44]
      reg_inst <= 32'h0; // @[PipelineReg.scala 39:14]
    end else if (_T) begin // @[PipelineReg.scala 86:27]
      reg_inst <= io_in_inst; // @[PipelineReg.scala 87:9]
    end
    if (reset) begin // @[PipelineReg.scala 82:20]
      reg_typeL <= 1'h0; // @[PipelineReg.scala 82:20]
    end else if (io_flush & ~io_stall) begin // @[PipelineReg.scala 84:44]
      reg_typeL <= 1'h0; // @[PipelineReg.scala 40:14]
    end else if (_T) begin // @[PipelineReg.scala 86:27]
      reg_typeL <= io_in_typeL; // @[PipelineReg.scala 87:9]
    end
    if (reset) begin // @[PipelineReg.scala 82:20]
      reg_aluA <= 1'h0; // @[PipelineReg.scala 82:20]
    end else if (io_flush & ~io_stall) begin // @[PipelineReg.scala 84:44]
      reg_aluA <= 1'h0; // @[PipelineReg.scala 42:14]
    end else if (_T) begin // @[PipelineReg.scala 86:27]
      reg_aluA <= io_in_aluA; // @[PipelineReg.scala 87:9]
    end
    if (reset) begin // @[PipelineReg.scala 82:20]
      reg_aluB <= 2'h0; // @[PipelineReg.scala 82:20]
    end else if (io_flush & ~io_stall) begin // @[PipelineReg.scala 84:44]
      reg_aluB <= 2'h3; // @[PipelineReg.scala 43:14]
    end else if (_T) begin // @[PipelineReg.scala 86:27]
      reg_aluB <= io_in_aluB; // @[PipelineReg.scala 87:9]
    end
    if (reset) begin // @[PipelineReg.scala 82:20]
      reg_aluOp <= 4'h0; // @[PipelineReg.scala 82:20]
    end else if (io_flush & ~io_stall) begin // @[PipelineReg.scala 84:44]
      reg_aluOp <= 4'h0; // @[PipelineReg.scala 44:14]
    end else if (_T) begin // @[PipelineReg.scala 86:27]
      reg_aluOp <= io_in_aluOp; // @[PipelineReg.scala 87:9]
    end
    if (reset) begin // @[PipelineReg.scala 82:20]
      reg_branch <= 3'h0; // @[PipelineReg.scala 82:20]
    end else if (io_flush & ~io_stall) begin // @[PipelineReg.scala 84:44]
      reg_branch <= 3'h0; // @[PipelineReg.scala 46:14]
    end else if (_T) begin // @[PipelineReg.scala 86:27]
      reg_branch <= io_in_branch; // @[PipelineReg.scala 87:9]
    end
    if (reset) begin // @[PipelineReg.scala 82:20]
      reg_memtoReg <= 2'h0; // @[PipelineReg.scala 82:20]
    end else if (io_flush & ~io_stall) begin // @[PipelineReg.scala 84:44]
      reg_memtoReg <= 2'h0; // @[PipelineReg.scala 47:14]
    end else if (_T) begin // @[PipelineReg.scala 86:27]
      reg_memtoReg <= io_in_memtoReg; // @[PipelineReg.scala 87:9]
    end
    if (reset) begin // @[PipelineReg.scala 82:20]
      reg_memWr <= 1'h0; // @[PipelineReg.scala 82:20]
    end else if (io_flush & ~io_stall) begin // @[PipelineReg.scala 84:44]
      reg_memWr <= 1'h0; // @[PipelineReg.scala 48:14]
    end else if (_T) begin // @[PipelineReg.scala 86:27]
      reg_memWr <= io_in_memWr; // @[PipelineReg.scala 87:9]
    end
    if (reset) begin // @[PipelineReg.scala 82:20]
      reg_memOp <= 3'h0; // @[PipelineReg.scala 82:20]
    end else if (io_flush & ~io_stall) begin // @[PipelineReg.scala 84:44]
      reg_memOp <= 3'h0; // @[PipelineReg.scala 49:14]
    end else if (_T) begin // @[PipelineReg.scala 86:27]
      reg_memOp <= io_in_memOp; // @[PipelineReg.scala 87:9]
    end
    if (reset) begin // @[PipelineReg.scala 82:20]
      reg_memAddr <= 32'h0; // @[PipelineReg.scala 82:20]
    end else if (io_flush & ~io_stall) begin // @[PipelineReg.scala 84:44]
      reg_memAddr <= 32'h0; // @[PipelineReg.scala 50:14]
    end else if (_T) begin // @[PipelineReg.scala 86:27]
      reg_memAddr <= io_in_memAddr; // @[PipelineReg.scala 87:9]
    end
    if (reset) begin // @[PipelineReg.scala 82:20]
      reg_rdEn <= 1'h0; // @[PipelineReg.scala 82:20]
    end else if (io_flush & ~io_stall) begin // @[PipelineReg.scala 84:44]
      reg_rdEn <= 1'h0; // @[PipelineReg.scala 52:14]
    end else if (_T) begin // @[PipelineReg.scala 86:27]
      reg_rdEn <= io_in_rdEn; // @[PipelineReg.scala 87:9]
    end
    if (reset) begin // @[PipelineReg.scala 82:20]
      reg_rdAddr <= 5'h0; // @[PipelineReg.scala 82:20]
    end else if (io_flush & ~io_stall) begin // @[PipelineReg.scala 84:44]
      reg_rdAddr <= 5'h0; // @[PipelineReg.scala 53:14]
    end else if (_T) begin // @[PipelineReg.scala 86:27]
      reg_rdAddr <= io_in_rdAddr; // @[PipelineReg.scala 87:9]
    end
    if (reset) begin // @[PipelineReg.scala 82:20]
      reg_rs1Data <= 64'h0; // @[PipelineReg.scala 82:20]
    end else if (io_flush & ~io_stall) begin // @[PipelineReg.scala 84:44]
      reg_rs1Data <= 64'h0; // @[PipelineReg.scala 54:14]
    end else if (_T) begin // @[PipelineReg.scala 86:27]
      reg_rs1Data <= io_in_rs1Data; // @[PipelineReg.scala 87:9]
    end
    if (reset) begin // @[PipelineReg.scala 82:20]
      reg_rs2Data <= 64'h0; // @[PipelineReg.scala 82:20]
    end else if (io_flush & ~io_stall) begin // @[PipelineReg.scala 84:44]
      reg_rs2Data <= 64'h0; // @[PipelineReg.scala 55:14]
    end else if (_T) begin // @[PipelineReg.scala 86:27]
      reg_rs2Data <= io_in_rs2Data; // @[PipelineReg.scala 87:9]
    end
    if (reset) begin // @[PipelineReg.scala 82:20]
      reg_imm <= 64'h0; // @[PipelineReg.scala 82:20]
    end else if (io_flush & ~io_stall) begin // @[PipelineReg.scala 84:44]
      reg_imm <= 64'h0; // @[PipelineReg.scala 56:14]
    end else if (_T) begin // @[PipelineReg.scala 86:27]
      reg_imm <= io_in_imm; // @[PipelineReg.scala 87:9]
    end
    if (reset) begin // @[PipelineReg.scala 82:20]
      reg_aluRes <= 64'h0; // @[PipelineReg.scala 82:20]
    end else if (io_flush & ~io_stall) begin // @[PipelineReg.scala 84:44]
      reg_aluRes <= 64'h0; // @[PipelineReg.scala 60:14]
    end else if (_T) begin // @[PipelineReg.scala 86:27]
      reg_aluRes <= io_in_aluRes; // @[PipelineReg.scala 87:9]
    end
    if (reset) begin // @[PipelineReg.scala 82:20]
      reg_memData <= 64'h0; // @[PipelineReg.scala 82:20]
    end else if (io_flush & ~io_stall) begin // @[PipelineReg.scala 84:44]
      reg_memData <= 64'h0; // @[PipelineReg.scala 61:14]
    end else if (_T) begin // @[PipelineReg.scala 86:27]
      reg_memData <= io_in_memData; // @[PipelineReg.scala 87:9]
    end
    if (reset) begin // @[PipelineReg.scala 82:20]
      reg_csrOp <= 4'h0; // @[PipelineReg.scala 82:20]
    end else if (io_flush & ~io_stall) begin // @[PipelineReg.scala 84:44]
      reg_csrOp <= 4'h0; // @[PipelineReg.scala 63:11]
    end else if (_T) begin // @[PipelineReg.scala 86:27]
      reg_csrOp <= io_in_csrOp; // @[PipelineReg.scala 87:9]
    end
    if (reset) begin // @[PipelineReg.scala 82:20]
      reg_takenPre <= 1'h0; // @[PipelineReg.scala 82:20]
    end else if (io_flush & ~io_stall) begin // @[PipelineReg.scala 84:44]
      reg_takenPre <= 1'h0; // @[PipelineReg.scala 65:15]
    end else if (_T) begin // @[PipelineReg.scala 86:27]
      reg_takenPre <= io_in_takenPre; // @[PipelineReg.scala 87:9]
    end
    if (reset) begin // @[PipelineReg.scala 82:20]
      reg_takenPrePC <= 32'h0; // @[PipelineReg.scala 82:20]
    end else if (io_flush & ~io_stall) begin // @[PipelineReg.scala 84:44]
      reg_takenPrePC <= 32'h0; // @[PipelineReg.scala 66:16]
    end else if (_T) begin // @[PipelineReg.scala 86:27]
      reg_takenPrePC <= io_in_takenPrePC; // @[PipelineReg.scala 87:9]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reg_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  reg_pc = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  reg_inst = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  reg_typeL = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  reg_aluA = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  reg_aluB = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  reg_aluOp = _RAND_6[3:0];
  _RAND_7 = {1{`RANDOM}};
  reg_branch = _RAND_7[2:0];
  _RAND_8 = {1{`RANDOM}};
  reg_memtoReg = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  reg_memWr = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  reg_memOp = _RAND_10[2:0];
  _RAND_11 = {1{`RANDOM}};
  reg_memAddr = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  reg_rdEn = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  reg_rdAddr = _RAND_13[4:0];
  _RAND_14 = {2{`RANDOM}};
  reg_rs1Data = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  reg_rs2Data = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  reg_imm = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  reg_aluRes = _RAND_17[63:0];
  _RAND_18 = {2{`RANDOM}};
  reg_memData = _RAND_18[63:0];
  _RAND_19 = {1{`RANDOM}};
  reg_csrOp = _RAND_19[3:0];
  _RAND_20 = {1{`RANDOM}};
  reg_takenPre = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  reg_takenPrePC = _RAND_21[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RegFile(
  input         clock,
  input         reset,
  output [63:0] io_rs1Data,
  output [63:0] io_rs2Data,
  input         io_rdEn,
  input  [31:0] io_rdAddr,
  input  [63:0] io_rdData,
  input         io_preRs1En,
  input  [4:0]  io_preRs1Addr,
  output [63:0] io_preRs1Data,
  output [63:0] io_preRs1x1Data,
  input         io_ctrl_rs1En,
  input         io_ctrl_rs2En,
  input  [4:0]  io_ctrl_rs1Addr,
  input  [4:0]  io_ctrl_rs2Addr,
  output [63:0] rf_10
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
`endif // RANDOMIZE_REG_INIT
  wire  dt_ar_clock; // @[RegFile.scala 36:21]
  wire [7:0] dt_ar_coreid; // @[RegFile.scala 36:21]
  wire [63:0] dt_ar_gpr_0; // @[RegFile.scala 36:21]
  wire [63:0] dt_ar_gpr_1; // @[RegFile.scala 36:21]
  wire [63:0] dt_ar_gpr_2; // @[RegFile.scala 36:21]
  wire [63:0] dt_ar_gpr_3; // @[RegFile.scala 36:21]
  wire [63:0] dt_ar_gpr_4; // @[RegFile.scala 36:21]
  wire [63:0] dt_ar_gpr_5; // @[RegFile.scala 36:21]
  wire [63:0] dt_ar_gpr_6; // @[RegFile.scala 36:21]
  wire [63:0] dt_ar_gpr_7; // @[RegFile.scala 36:21]
  wire [63:0] dt_ar_gpr_8; // @[RegFile.scala 36:21]
  wire [63:0] dt_ar_gpr_9; // @[RegFile.scala 36:21]
  wire [63:0] dt_ar_gpr_10; // @[RegFile.scala 36:21]
  wire [63:0] dt_ar_gpr_11; // @[RegFile.scala 36:21]
  wire [63:0] dt_ar_gpr_12; // @[RegFile.scala 36:21]
  wire [63:0] dt_ar_gpr_13; // @[RegFile.scala 36:21]
  wire [63:0] dt_ar_gpr_14; // @[RegFile.scala 36:21]
  wire [63:0] dt_ar_gpr_15; // @[RegFile.scala 36:21]
  wire [63:0] dt_ar_gpr_16; // @[RegFile.scala 36:21]
  wire [63:0] dt_ar_gpr_17; // @[RegFile.scala 36:21]
  wire [63:0] dt_ar_gpr_18; // @[RegFile.scala 36:21]
  wire [63:0] dt_ar_gpr_19; // @[RegFile.scala 36:21]
  wire [63:0] dt_ar_gpr_20; // @[RegFile.scala 36:21]
  wire [63:0] dt_ar_gpr_21; // @[RegFile.scala 36:21]
  wire [63:0] dt_ar_gpr_22; // @[RegFile.scala 36:21]
  wire [63:0] dt_ar_gpr_23; // @[RegFile.scala 36:21]
  wire [63:0] dt_ar_gpr_24; // @[RegFile.scala 36:21]
  wire [63:0] dt_ar_gpr_25; // @[RegFile.scala 36:21]
  wire [63:0] dt_ar_gpr_26; // @[RegFile.scala 36:21]
  wire [63:0] dt_ar_gpr_27; // @[RegFile.scala 36:21]
  wire [63:0] dt_ar_gpr_28; // @[RegFile.scala 36:21]
  wire [63:0] dt_ar_gpr_29; // @[RegFile.scala 36:21]
  wire [63:0] dt_ar_gpr_30; // @[RegFile.scala 36:21]
  wire [63:0] dt_ar_gpr_31; // @[RegFile.scala 36:21]
  reg [63:0] rf__0; // @[RegFile.scala 24:19]
  reg [63:0] rf__1; // @[RegFile.scala 24:19]
  reg [63:0] rf__2; // @[RegFile.scala 24:19]
  reg [63:0] rf__3; // @[RegFile.scala 24:19]
  reg [63:0] rf__4; // @[RegFile.scala 24:19]
  reg [63:0] rf__5; // @[RegFile.scala 24:19]
  reg [63:0] rf__6; // @[RegFile.scala 24:19]
  reg [63:0] rf__7; // @[RegFile.scala 24:19]
  reg [63:0] rf__8; // @[RegFile.scala 24:19]
  reg [63:0] rf__9; // @[RegFile.scala 24:19]
  reg [63:0] rf__10; // @[RegFile.scala 24:19]
  reg [63:0] rf__11; // @[RegFile.scala 24:19]
  reg [63:0] rf__12; // @[RegFile.scala 24:19]
  reg [63:0] rf__13; // @[RegFile.scala 24:19]
  reg [63:0] rf__14; // @[RegFile.scala 24:19]
  reg [63:0] rf__15; // @[RegFile.scala 24:19]
  reg [63:0] rf__16; // @[RegFile.scala 24:19]
  reg [63:0] rf__17; // @[RegFile.scala 24:19]
  reg [63:0] rf__18; // @[RegFile.scala 24:19]
  reg [63:0] rf__19; // @[RegFile.scala 24:19]
  reg [63:0] rf__20; // @[RegFile.scala 24:19]
  reg [63:0] rf__21; // @[RegFile.scala 24:19]
  reg [63:0] rf__22; // @[RegFile.scala 24:19]
  reg [63:0] rf__23; // @[RegFile.scala 24:19]
  reg [63:0] rf__24; // @[RegFile.scala 24:19]
  reg [63:0] rf__25; // @[RegFile.scala 24:19]
  reg [63:0] rf__26; // @[RegFile.scala 24:19]
  reg [63:0] rf__27; // @[RegFile.scala 24:19]
  reg [63:0] rf__28; // @[RegFile.scala 24:19]
  reg [63:0] rf__29; // @[RegFile.scala 24:19]
  reg [63:0] rf__30; // @[RegFile.scala 24:19]
  reg [63:0] rf__31; // @[RegFile.scala 24:19]
  wire [63:0] _GEN_65 = 5'h1 == io_ctrl_rs1Addr ? rf__1 : rf__0; // @[RegFile.scala 30:{20,20}]
  wire [63:0] _GEN_66 = 5'h2 == io_ctrl_rs1Addr ? rf__2 : _GEN_65; // @[RegFile.scala 30:{20,20}]
  wire [63:0] _GEN_67 = 5'h3 == io_ctrl_rs1Addr ? rf__3 : _GEN_66; // @[RegFile.scala 30:{20,20}]
  wire [63:0] _GEN_68 = 5'h4 == io_ctrl_rs1Addr ? rf__4 : _GEN_67; // @[RegFile.scala 30:{20,20}]
  wire [63:0] _GEN_69 = 5'h5 == io_ctrl_rs1Addr ? rf__5 : _GEN_68; // @[RegFile.scala 30:{20,20}]
  wire [63:0] _GEN_70 = 5'h6 == io_ctrl_rs1Addr ? rf__6 : _GEN_69; // @[RegFile.scala 30:{20,20}]
  wire [63:0] _GEN_71 = 5'h7 == io_ctrl_rs1Addr ? rf__7 : _GEN_70; // @[RegFile.scala 30:{20,20}]
  wire [63:0] _GEN_72 = 5'h8 == io_ctrl_rs1Addr ? rf__8 : _GEN_71; // @[RegFile.scala 30:{20,20}]
  wire [63:0] _GEN_73 = 5'h9 == io_ctrl_rs1Addr ? rf__9 : _GEN_72; // @[RegFile.scala 30:{20,20}]
  wire [63:0] _GEN_74 = 5'ha == io_ctrl_rs1Addr ? rf__10 : _GEN_73; // @[RegFile.scala 30:{20,20}]
  wire [63:0] _GEN_75 = 5'hb == io_ctrl_rs1Addr ? rf__11 : _GEN_74; // @[RegFile.scala 30:{20,20}]
  wire [63:0] _GEN_76 = 5'hc == io_ctrl_rs1Addr ? rf__12 : _GEN_75; // @[RegFile.scala 30:{20,20}]
  wire [63:0] _GEN_77 = 5'hd == io_ctrl_rs1Addr ? rf__13 : _GEN_76; // @[RegFile.scala 30:{20,20}]
  wire [63:0] _GEN_78 = 5'he == io_ctrl_rs1Addr ? rf__14 : _GEN_77; // @[RegFile.scala 30:{20,20}]
  wire [63:0] _GEN_79 = 5'hf == io_ctrl_rs1Addr ? rf__15 : _GEN_78; // @[RegFile.scala 30:{20,20}]
  wire [63:0] _GEN_80 = 5'h10 == io_ctrl_rs1Addr ? rf__16 : _GEN_79; // @[RegFile.scala 30:{20,20}]
  wire [63:0] _GEN_81 = 5'h11 == io_ctrl_rs1Addr ? rf__17 : _GEN_80; // @[RegFile.scala 30:{20,20}]
  wire [63:0] _GEN_82 = 5'h12 == io_ctrl_rs1Addr ? rf__18 : _GEN_81; // @[RegFile.scala 30:{20,20}]
  wire [63:0] _GEN_83 = 5'h13 == io_ctrl_rs1Addr ? rf__19 : _GEN_82; // @[RegFile.scala 30:{20,20}]
  wire [63:0] _GEN_84 = 5'h14 == io_ctrl_rs1Addr ? rf__20 : _GEN_83; // @[RegFile.scala 30:{20,20}]
  wire [63:0] _GEN_85 = 5'h15 == io_ctrl_rs1Addr ? rf__21 : _GEN_84; // @[RegFile.scala 30:{20,20}]
  wire [63:0] _GEN_86 = 5'h16 == io_ctrl_rs1Addr ? rf__22 : _GEN_85; // @[RegFile.scala 30:{20,20}]
  wire [63:0] _GEN_87 = 5'h17 == io_ctrl_rs1Addr ? rf__23 : _GEN_86; // @[RegFile.scala 30:{20,20}]
  wire [63:0] _GEN_88 = 5'h18 == io_ctrl_rs1Addr ? rf__24 : _GEN_87; // @[RegFile.scala 30:{20,20}]
  wire [63:0] _GEN_89 = 5'h19 == io_ctrl_rs1Addr ? rf__25 : _GEN_88; // @[RegFile.scala 30:{20,20}]
  wire [63:0] _GEN_90 = 5'h1a == io_ctrl_rs1Addr ? rf__26 : _GEN_89; // @[RegFile.scala 30:{20,20}]
  wire [63:0] _GEN_91 = 5'h1b == io_ctrl_rs1Addr ? rf__27 : _GEN_90; // @[RegFile.scala 30:{20,20}]
  wire [63:0] _GEN_92 = 5'h1c == io_ctrl_rs1Addr ? rf__28 : _GEN_91; // @[RegFile.scala 30:{20,20}]
  wire [63:0] _GEN_93 = 5'h1d == io_ctrl_rs1Addr ? rf__29 : _GEN_92; // @[RegFile.scala 30:{20,20}]
  wire [63:0] _GEN_94 = 5'h1e == io_ctrl_rs1Addr ? rf__30 : _GEN_93; // @[RegFile.scala 30:{20,20}]
  wire [63:0] _GEN_95 = 5'h1f == io_ctrl_rs1Addr ? rf__31 : _GEN_94; // @[RegFile.scala 30:{20,20}]
  wire [63:0] _GEN_97 = 5'h1 == io_ctrl_rs2Addr ? rf__1 : rf__0; // @[RegFile.scala 31:{20,20}]
  wire [63:0] _GEN_98 = 5'h2 == io_ctrl_rs2Addr ? rf__2 : _GEN_97; // @[RegFile.scala 31:{20,20}]
  wire [63:0] _GEN_99 = 5'h3 == io_ctrl_rs2Addr ? rf__3 : _GEN_98; // @[RegFile.scala 31:{20,20}]
  wire [63:0] _GEN_100 = 5'h4 == io_ctrl_rs2Addr ? rf__4 : _GEN_99; // @[RegFile.scala 31:{20,20}]
  wire [63:0] _GEN_101 = 5'h5 == io_ctrl_rs2Addr ? rf__5 : _GEN_100; // @[RegFile.scala 31:{20,20}]
  wire [63:0] _GEN_102 = 5'h6 == io_ctrl_rs2Addr ? rf__6 : _GEN_101; // @[RegFile.scala 31:{20,20}]
  wire [63:0] _GEN_103 = 5'h7 == io_ctrl_rs2Addr ? rf__7 : _GEN_102; // @[RegFile.scala 31:{20,20}]
  wire [63:0] _GEN_104 = 5'h8 == io_ctrl_rs2Addr ? rf__8 : _GEN_103; // @[RegFile.scala 31:{20,20}]
  wire [63:0] _GEN_105 = 5'h9 == io_ctrl_rs2Addr ? rf__9 : _GEN_104; // @[RegFile.scala 31:{20,20}]
  wire [63:0] _GEN_106 = 5'ha == io_ctrl_rs2Addr ? rf__10 : _GEN_105; // @[RegFile.scala 31:{20,20}]
  wire [63:0] _GEN_107 = 5'hb == io_ctrl_rs2Addr ? rf__11 : _GEN_106; // @[RegFile.scala 31:{20,20}]
  wire [63:0] _GEN_108 = 5'hc == io_ctrl_rs2Addr ? rf__12 : _GEN_107; // @[RegFile.scala 31:{20,20}]
  wire [63:0] _GEN_109 = 5'hd == io_ctrl_rs2Addr ? rf__13 : _GEN_108; // @[RegFile.scala 31:{20,20}]
  wire [63:0] _GEN_110 = 5'he == io_ctrl_rs2Addr ? rf__14 : _GEN_109; // @[RegFile.scala 31:{20,20}]
  wire [63:0] _GEN_111 = 5'hf == io_ctrl_rs2Addr ? rf__15 : _GEN_110; // @[RegFile.scala 31:{20,20}]
  wire [63:0] _GEN_112 = 5'h10 == io_ctrl_rs2Addr ? rf__16 : _GEN_111; // @[RegFile.scala 31:{20,20}]
  wire [63:0] _GEN_113 = 5'h11 == io_ctrl_rs2Addr ? rf__17 : _GEN_112; // @[RegFile.scala 31:{20,20}]
  wire [63:0] _GEN_114 = 5'h12 == io_ctrl_rs2Addr ? rf__18 : _GEN_113; // @[RegFile.scala 31:{20,20}]
  wire [63:0] _GEN_115 = 5'h13 == io_ctrl_rs2Addr ? rf__19 : _GEN_114; // @[RegFile.scala 31:{20,20}]
  wire [63:0] _GEN_116 = 5'h14 == io_ctrl_rs2Addr ? rf__20 : _GEN_115; // @[RegFile.scala 31:{20,20}]
  wire [63:0] _GEN_117 = 5'h15 == io_ctrl_rs2Addr ? rf__21 : _GEN_116; // @[RegFile.scala 31:{20,20}]
  wire [63:0] _GEN_118 = 5'h16 == io_ctrl_rs2Addr ? rf__22 : _GEN_117; // @[RegFile.scala 31:{20,20}]
  wire [63:0] _GEN_119 = 5'h17 == io_ctrl_rs2Addr ? rf__23 : _GEN_118; // @[RegFile.scala 31:{20,20}]
  wire [63:0] _GEN_120 = 5'h18 == io_ctrl_rs2Addr ? rf__24 : _GEN_119; // @[RegFile.scala 31:{20,20}]
  wire [63:0] _GEN_121 = 5'h19 == io_ctrl_rs2Addr ? rf__25 : _GEN_120; // @[RegFile.scala 31:{20,20}]
  wire [63:0] _GEN_122 = 5'h1a == io_ctrl_rs2Addr ? rf__26 : _GEN_121; // @[RegFile.scala 31:{20,20}]
  wire [63:0] _GEN_123 = 5'h1b == io_ctrl_rs2Addr ? rf__27 : _GEN_122; // @[RegFile.scala 31:{20,20}]
  wire [63:0] _GEN_124 = 5'h1c == io_ctrl_rs2Addr ? rf__28 : _GEN_123; // @[RegFile.scala 31:{20,20}]
  wire [63:0] _GEN_125 = 5'h1d == io_ctrl_rs2Addr ? rf__29 : _GEN_124; // @[RegFile.scala 31:{20,20}]
  wire [63:0] _GEN_126 = 5'h1e == io_ctrl_rs2Addr ? rf__30 : _GEN_125; // @[RegFile.scala 31:{20,20}]
  wire [63:0] _GEN_127 = 5'h1f == io_ctrl_rs2Addr ? rf__31 : _GEN_126; // @[RegFile.scala 31:{20,20}]
  wire [63:0] _GEN_129 = 5'h1 == io_preRs1Addr ? rf__1 : rf__0; // @[RegFile.scala 34:{23,23}]
  wire [63:0] _GEN_130 = 5'h2 == io_preRs1Addr ? rf__2 : _GEN_129; // @[RegFile.scala 34:{23,23}]
  wire [63:0] _GEN_131 = 5'h3 == io_preRs1Addr ? rf__3 : _GEN_130; // @[RegFile.scala 34:{23,23}]
  wire [63:0] _GEN_132 = 5'h4 == io_preRs1Addr ? rf__4 : _GEN_131; // @[RegFile.scala 34:{23,23}]
  wire [63:0] _GEN_133 = 5'h5 == io_preRs1Addr ? rf__5 : _GEN_132; // @[RegFile.scala 34:{23,23}]
  wire [63:0] _GEN_134 = 5'h6 == io_preRs1Addr ? rf__6 : _GEN_133; // @[RegFile.scala 34:{23,23}]
  wire [63:0] _GEN_135 = 5'h7 == io_preRs1Addr ? rf__7 : _GEN_134; // @[RegFile.scala 34:{23,23}]
  wire [63:0] _GEN_136 = 5'h8 == io_preRs1Addr ? rf__8 : _GEN_135; // @[RegFile.scala 34:{23,23}]
  wire [63:0] _GEN_137 = 5'h9 == io_preRs1Addr ? rf__9 : _GEN_136; // @[RegFile.scala 34:{23,23}]
  wire [63:0] _GEN_138 = 5'ha == io_preRs1Addr ? rf__10 : _GEN_137; // @[RegFile.scala 34:{23,23}]
  wire [63:0] _GEN_139 = 5'hb == io_preRs1Addr ? rf__11 : _GEN_138; // @[RegFile.scala 34:{23,23}]
  wire [63:0] _GEN_140 = 5'hc == io_preRs1Addr ? rf__12 : _GEN_139; // @[RegFile.scala 34:{23,23}]
  wire [63:0] _GEN_141 = 5'hd == io_preRs1Addr ? rf__13 : _GEN_140; // @[RegFile.scala 34:{23,23}]
  wire [63:0] _GEN_142 = 5'he == io_preRs1Addr ? rf__14 : _GEN_141; // @[RegFile.scala 34:{23,23}]
  wire [63:0] _GEN_143 = 5'hf == io_preRs1Addr ? rf__15 : _GEN_142; // @[RegFile.scala 34:{23,23}]
  wire [63:0] _GEN_144 = 5'h10 == io_preRs1Addr ? rf__16 : _GEN_143; // @[RegFile.scala 34:{23,23}]
  wire [63:0] _GEN_145 = 5'h11 == io_preRs1Addr ? rf__17 : _GEN_144; // @[RegFile.scala 34:{23,23}]
  wire [63:0] _GEN_146 = 5'h12 == io_preRs1Addr ? rf__18 : _GEN_145; // @[RegFile.scala 34:{23,23}]
  wire [63:0] _GEN_147 = 5'h13 == io_preRs1Addr ? rf__19 : _GEN_146; // @[RegFile.scala 34:{23,23}]
  wire [63:0] _GEN_148 = 5'h14 == io_preRs1Addr ? rf__20 : _GEN_147; // @[RegFile.scala 34:{23,23}]
  wire [63:0] _GEN_149 = 5'h15 == io_preRs1Addr ? rf__21 : _GEN_148; // @[RegFile.scala 34:{23,23}]
  wire [63:0] _GEN_150 = 5'h16 == io_preRs1Addr ? rf__22 : _GEN_149; // @[RegFile.scala 34:{23,23}]
  wire [63:0] _GEN_151 = 5'h17 == io_preRs1Addr ? rf__23 : _GEN_150; // @[RegFile.scala 34:{23,23}]
  wire [63:0] _GEN_152 = 5'h18 == io_preRs1Addr ? rf__24 : _GEN_151; // @[RegFile.scala 34:{23,23}]
  wire [63:0] _GEN_153 = 5'h19 == io_preRs1Addr ? rf__25 : _GEN_152; // @[RegFile.scala 34:{23,23}]
  wire [63:0] _GEN_154 = 5'h1a == io_preRs1Addr ? rf__26 : _GEN_153; // @[RegFile.scala 34:{23,23}]
  wire [63:0] _GEN_155 = 5'h1b == io_preRs1Addr ? rf__27 : _GEN_154; // @[RegFile.scala 34:{23,23}]
  wire [63:0] _GEN_156 = 5'h1c == io_preRs1Addr ? rf__28 : _GEN_155; // @[RegFile.scala 34:{23,23}]
  wire [63:0] _GEN_157 = 5'h1d == io_preRs1Addr ? rf__29 : _GEN_156; // @[RegFile.scala 34:{23,23}]
  wire [63:0] _GEN_158 = 5'h1e == io_preRs1Addr ? rf__30 : _GEN_157; // @[RegFile.scala 34:{23,23}]
  wire [63:0] _GEN_159 = 5'h1f == io_preRs1Addr ? rf__31 : _GEN_158; // @[RegFile.scala 34:{23,23}]
  DifftestArchIntRegState dt_ar ( // @[RegFile.scala 36:21]
    .clock(dt_ar_clock),
    .coreid(dt_ar_coreid),
    .gpr_0(dt_ar_gpr_0),
    .gpr_1(dt_ar_gpr_1),
    .gpr_2(dt_ar_gpr_2),
    .gpr_3(dt_ar_gpr_3),
    .gpr_4(dt_ar_gpr_4),
    .gpr_5(dt_ar_gpr_5),
    .gpr_6(dt_ar_gpr_6),
    .gpr_7(dt_ar_gpr_7),
    .gpr_8(dt_ar_gpr_8),
    .gpr_9(dt_ar_gpr_9),
    .gpr_10(dt_ar_gpr_10),
    .gpr_11(dt_ar_gpr_11),
    .gpr_12(dt_ar_gpr_12),
    .gpr_13(dt_ar_gpr_13),
    .gpr_14(dt_ar_gpr_14),
    .gpr_15(dt_ar_gpr_15),
    .gpr_16(dt_ar_gpr_16),
    .gpr_17(dt_ar_gpr_17),
    .gpr_18(dt_ar_gpr_18),
    .gpr_19(dt_ar_gpr_19),
    .gpr_20(dt_ar_gpr_20),
    .gpr_21(dt_ar_gpr_21),
    .gpr_22(dt_ar_gpr_22),
    .gpr_23(dt_ar_gpr_23),
    .gpr_24(dt_ar_gpr_24),
    .gpr_25(dt_ar_gpr_25),
    .gpr_26(dt_ar_gpr_26),
    .gpr_27(dt_ar_gpr_27),
    .gpr_28(dt_ar_gpr_28),
    .gpr_29(dt_ar_gpr_29),
    .gpr_30(dt_ar_gpr_30),
    .gpr_31(dt_ar_gpr_31)
  );
  assign io_rs1Data = io_ctrl_rs1Addr != 5'h0 & io_ctrl_rs1En ? _GEN_95 : 64'h0; // @[RegFile.scala 30:20]
  assign io_rs2Data = io_ctrl_rs2Addr != 5'h0 & io_ctrl_rs2En ? _GEN_127 : 64'h0; // @[RegFile.scala 31:20]
  assign io_preRs1Data = io_preRs1En & io_preRs1Addr != 5'h0 & io_preRs1Addr != 5'h1 ? _GEN_159 : 64'h0; // @[RegFile.scala 34:23]
  assign io_preRs1x1Data = rf__1; // @[RegFile.scala 33:19]
  assign rf_10 = rf__10;
  assign dt_ar_clock = clock; // @[RegFile.scala 37:19]
  assign dt_ar_coreid = 8'h0; // @[RegFile.scala 38:19]
  assign dt_ar_gpr_0 = rf__0; // @[RegFile.scala 39:19]
  assign dt_ar_gpr_1 = rf__1; // @[RegFile.scala 39:19]
  assign dt_ar_gpr_2 = rf__2; // @[RegFile.scala 39:19]
  assign dt_ar_gpr_3 = rf__3; // @[RegFile.scala 39:19]
  assign dt_ar_gpr_4 = rf__4; // @[RegFile.scala 39:19]
  assign dt_ar_gpr_5 = rf__5; // @[RegFile.scala 39:19]
  assign dt_ar_gpr_6 = rf__6; // @[RegFile.scala 39:19]
  assign dt_ar_gpr_7 = rf__7; // @[RegFile.scala 39:19]
  assign dt_ar_gpr_8 = rf__8; // @[RegFile.scala 39:19]
  assign dt_ar_gpr_9 = rf__9; // @[RegFile.scala 39:19]
  assign dt_ar_gpr_10 = rf__10; // @[RegFile.scala 39:19]
  assign dt_ar_gpr_11 = rf__11; // @[RegFile.scala 39:19]
  assign dt_ar_gpr_12 = rf__12; // @[RegFile.scala 39:19]
  assign dt_ar_gpr_13 = rf__13; // @[RegFile.scala 39:19]
  assign dt_ar_gpr_14 = rf__14; // @[RegFile.scala 39:19]
  assign dt_ar_gpr_15 = rf__15; // @[RegFile.scala 39:19]
  assign dt_ar_gpr_16 = rf__16; // @[RegFile.scala 39:19]
  assign dt_ar_gpr_17 = rf__17; // @[RegFile.scala 39:19]
  assign dt_ar_gpr_18 = rf__18; // @[RegFile.scala 39:19]
  assign dt_ar_gpr_19 = rf__19; // @[RegFile.scala 39:19]
  assign dt_ar_gpr_20 = rf__20; // @[RegFile.scala 39:19]
  assign dt_ar_gpr_21 = rf__21; // @[RegFile.scala 39:19]
  assign dt_ar_gpr_22 = rf__22; // @[RegFile.scala 39:19]
  assign dt_ar_gpr_23 = rf__23; // @[RegFile.scala 39:19]
  assign dt_ar_gpr_24 = rf__24; // @[RegFile.scala 39:19]
  assign dt_ar_gpr_25 = rf__25; // @[RegFile.scala 39:19]
  assign dt_ar_gpr_26 = rf__26; // @[RegFile.scala 39:19]
  assign dt_ar_gpr_27 = rf__27; // @[RegFile.scala 39:19]
  assign dt_ar_gpr_28 = rf__28; // @[RegFile.scala 39:19]
  assign dt_ar_gpr_29 = rf__29; // @[RegFile.scala 39:19]
  assign dt_ar_gpr_30 = rf__30; // @[RegFile.scala 39:19]
  assign dt_ar_gpr_31 = rf__31; // @[RegFile.scala 39:19]
  always @(posedge clock) begin
    if (reset) begin // @[RegFile.scala 24:19]
      rf__0 <= 64'h0; // @[RegFile.scala 24:19]
    end else if (io_rdEn & io_rdAddr != 32'h0) begin // @[RegFile.scala 26:41]
      if (5'h0 == io_rdAddr[4:0]) begin // @[RegFile.scala 27:19]
        rf__0 <= io_rdData; // @[RegFile.scala 27:19]
      end
    end
    if (reset) begin // @[RegFile.scala 24:19]
      rf__1 <= 64'h0; // @[RegFile.scala 24:19]
    end else if (io_rdEn & io_rdAddr != 32'h0) begin // @[RegFile.scala 26:41]
      if (5'h1 == io_rdAddr[4:0]) begin // @[RegFile.scala 27:19]
        rf__1 <= io_rdData; // @[RegFile.scala 27:19]
      end
    end
    if (reset) begin // @[RegFile.scala 24:19]
      rf__2 <= 64'h0; // @[RegFile.scala 24:19]
    end else if (io_rdEn & io_rdAddr != 32'h0) begin // @[RegFile.scala 26:41]
      if (5'h2 == io_rdAddr[4:0]) begin // @[RegFile.scala 27:19]
        rf__2 <= io_rdData; // @[RegFile.scala 27:19]
      end
    end
    if (reset) begin // @[RegFile.scala 24:19]
      rf__3 <= 64'h0; // @[RegFile.scala 24:19]
    end else if (io_rdEn & io_rdAddr != 32'h0) begin // @[RegFile.scala 26:41]
      if (5'h3 == io_rdAddr[4:0]) begin // @[RegFile.scala 27:19]
        rf__3 <= io_rdData; // @[RegFile.scala 27:19]
      end
    end
    if (reset) begin // @[RegFile.scala 24:19]
      rf__4 <= 64'h0; // @[RegFile.scala 24:19]
    end else if (io_rdEn & io_rdAddr != 32'h0) begin // @[RegFile.scala 26:41]
      if (5'h4 == io_rdAddr[4:0]) begin // @[RegFile.scala 27:19]
        rf__4 <= io_rdData; // @[RegFile.scala 27:19]
      end
    end
    if (reset) begin // @[RegFile.scala 24:19]
      rf__5 <= 64'h0; // @[RegFile.scala 24:19]
    end else if (io_rdEn & io_rdAddr != 32'h0) begin // @[RegFile.scala 26:41]
      if (5'h5 == io_rdAddr[4:0]) begin // @[RegFile.scala 27:19]
        rf__5 <= io_rdData; // @[RegFile.scala 27:19]
      end
    end
    if (reset) begin // @[RegFile.scala 24:19]
      rf__6 <= 64'h0; // @[RegFile.scala 24:19]
    end else if (io_rdEn & io_rdAddr != 32'h0) begin // @[RegFile.scala 26:41]
      if (5'h6 == io_rdAddr[4:0]) begin // @[RegFile.scala 27:19]
        rf__6 <= io_rdData; // @[RegFile.scala 27:19]
      end
    end
    if (reset) begin // @[RegFile.scala 24:19]
      rf__7 <= 64'h0; // @[RegFile.scala 24:19]
    end else if (io_rdEn & io_rdAddr != 32'h0) begin // @[RegFile.scala 26:41]
      if (5'h7 == io_rdAddr[4:0]) begin // @[RegFile.scala 27:19]
        rf__7 <= io_rdData; // @[RegFile.scala 27:19]
      end
    end
    if (reset) begin // @[RegFile.scala 24:19]
      rf__8 <= 64'h0; // @[RegFile.scala 24:19]
    end else if (io_rdEn & io_rdAddr != 32'h0) begin // @[RegFile.scala 26:41]
      if (5'h8 == io_rdAddr[4:0]) begin // @[RegFile.scala 27:19]
        rf__8 <= io_rdData; // @[RegFile.scala 27:19]
      end
    end
    if (reset) begin // @[RegFile.scala 24:19]
      rf__9 <= 64'h0; // @[RegFile.scala 24:19]
    end else if (io_rdEn & io_rdAddr != 32'h0) begin // @[RegFile.scala 26:41]
      if (5'h9 == io_rdAddr[4:0]) begin // @[RegFile.scala 27:19]
        rf__9 <= io_rdData; // @[RegFile.scala 27:19]
      end
    end
    if (reset) begin // @[RegFile.scala 24:19]
      rf__10 <= 64'h0; // @[RegFile.scala 24:19]
    end else if (io_rdEn & io_rdAddr != 32'h0) begin // @[RegFile.scala 26:41]
      if (5'ha == io_rdAddr[4:0]) begin // @[RegFile.scala 27:19]
        rf__10 <= io_rdData; // @[RegFile.scala 27:19]
      end
    end
    if (reset) begin // @[RegFile.scala 24:19]
      rf__11 <= 64'h0; // @[RegFile.scala 24:19]
    end else if (io_rdEn & io_rdAddr != 32'h0) begin // @[RegFile.scala 26:41]
      if (5'hb == io_rdAddr[4:0]) begin // @[RegFile.scala 27:19]
        rf__11 <= io_rdData; // @[RegFile.scala 27:19]
      end
    end
    if (reset) begin // @[RegFile.scala 24:19]
      rf__12 <= 64'h0; // @[RegFile.scala 24:19]
    end else if (io_rdEn & io_rdAddr != 32'h0) begin // @[RegFile.scala 26:41]
      if (5'hc == io_rdAddr[4:0]) begin // @[RegFile.scala 27:19]
        rf__12 <= io_rdData; // @[RegFile.scala 27:19]
      end
    end
    if (reset) begin // @[RegFile.scala 24:19]
      rf__13 <= 64'h0; // @[RegFile.scala 24:19]
    end else if (io_rdEn & io_rdAddr != 32'h0) begin // @[RegFile.scala 26:41]
      if (5'hd == io_rdAddr[4:0]) begin // @[RegFile.scala 27:19]
        rf__13 <= io_rdData; // @[RegFile.scala 27:19]
      end
    end
    if (reset) begin // @[RegFile.scala 24:19]
      rf__14 <= 64'h0; // @[RegFile.scala 24:19]
    end else if (io_rdEn & io_rdAddr != 32'h0) begin // @[RegFile.scala 26:41]
      if (5'he == io_rdAddr[4:0]) begin // @[RegFile.scala 27:19]
        rf__14 <= io_rdData; // @[RegFile.scala 27:19]
      end
    end
    if (reset) begin // @[RegFile.scala 24:19]
      rf__15 <= 64'h0; // @[RegFile.scala 24:19]
    end else if (io_rdEn & io_rdAddr != 32'h0) begin // @[RegFile.scala 26:41]
      if (5'hf == io_rdAddr[4:0]) begin // @[RegFile.scala 27:19]
        rf__15 <= io_rdData; // @[RegFile.scala 27:19]
      end
    end
    if (reset) begin // @[RegFile.scala 24:19]
      rf__16 <= 64'h0; // @[RegFile.scala 24:19]
    end else if (io_rdEn & io_rdAddr != 32'h0) begin // @[RegFile.scala 26:41]
      if (5'h10 == io_rdAddr[4:0]) begin // @[RegFile.scala 27:19]
        rf__16 <= io_rdData; // @[RegFile.scala 27:19]
      end
    end
    if (reset) begin // @[RegFile.scala 24:19]
      rf__17 <= 64'h0; // @[RegFile.scala 24:19]
    end else if (io_rdEn & io_rdAddr != 32'h0) begin // @[RegFile.scala 26:41]
      if (5'h11 == io_rdAddr[4:0]) begin // @[RegFile.scala 27:19]
        rf__17 <= io_rdData; // @[RegFile.scala 27:19]
      end
    end
    if (reset) begin // @[RegFile.scala 24:19]
      rf__18 <= 64'h0; // @[RegFile.scala 24:19]
    end else if (io_rdEn & io_rdAddr != 32'h0) begin // @[RegFile.scala 26:41]
      if (5'h12 == io_rdAddr[4:0]) begin // @[RegFile.scala 27:19]
        rf__18 <= io_rdData; // @[RegFile.scala 27:19]
      end
    end
    if (reset) begin // @[RegFile.scala 24:19]
      rf__19 <= 64'h0; // @[RegFile.scala 24:19]
    end else if (io_rdEn & io_rdAddr != 32'h0) begin // @[RegFile.scala 26:41]
      if (5'h13 == io_rdAddr[4:0]) begin // @[RegFile.scala 27:19]
        rf__19 <= io_rdData; // @[RegFile.scala 27:19]
      end
    end
    if (reset) begin // @[RegFile.scala 24:19]
      rf__20 <= 64'h0; // @[RegFile.scala 24:19]
    end else if (io_rdEn & io_rdAddr != 32'h0) begin // @[RegFile.scala 26:41]
      if (5'h14 == io_rdAddr[4:0]) begin // @[RegFile.scala 27:19]
        rf__20 <= io_rdData; // @[RegFile.scala 27:19]
      end
    end
    if (reset) begin // @[RegFile.scala 24:19]
      rf__21 <= 64'h0; // @[RegFile.scala 24:19]
    end else if (io_rdEn & io_rdAddr != 32'h0) begin // @[RegFile.scala 26:41]
      if (5'h15 == io_rdAddr[4:0]) begin // @[RegFile.scala 27:19]
        rf__21 <= io_rdData; // @[RegFile.scala 27:19]
      end
    end
    if (reset) begin // @[RegFile.scala 24:19]
      rf__22 <= 64'h0; // @[RegFile.scala 24:19]
    end else if (io_rdEn & io_rdAddr != 32'h0) begin // @[RegFile.scala 26:41]
      if (5'h16 == io_rdAddr[4:0]) begin // @[RegFile.scala 27:19]
        rf__22 <= io_rdData; // @[RegFile.scala 27:19]
      end
    end
    if (reset) begin // @[RegFile.scala 24:19]
      rf__23 <= 64'h0; // @[RegFile.scala 24:19]
    end else if (io_rdEn & io_rdAddr != 32'h0) begin // @[RegFile.scala 26:41]
      if (5'h17 == io_rdAddr[4:0]) begin // @[RegFile.scala 27:19]
        rf__23 <= io_rdData; // @[RegFile.scala 27:19]
      end
    end
    if (reset) begin // @[RegFile.scala 24:19]
      rf__24 <= 64'h0; // @[RegFile.scala 24:19]
    end else if (io_rdEn & io_rdAddr != 32'h0) begin // @[RegFile.scala 26:41]
      if (5'h18 == io_rdAddr[4:0]) begin // @[RegFile.scala 27:19]
        rf__24 <= io_rdData; // @[RegFile.scala 27:19]
      end
    end
    if (reset) begin // @[RegFile.scala 24:19]
      rf__25 <= 64'h0; // @[RegFile.scala 24:19]
    end else if (io_rdEn & io_rdAddr != 32'h0) begin // @[RegFile.scala 26:41]
      if (5'h19 == io_rdAddr[4:0]) begin // @[RegFile.scala 27:19]
        rf__25 <= io_rdData; // @[RegFile.scala 27:19]
      end
    end
    if (reset) begin // @[RegFile.scala 24:19]
      rf__26 <= 64'h0; // @[RegFile.scala 24:19]
    end else if (io_rdEn & io_rdAddr != 32'h0) begin // @[RegFile.scala 26:41]
      if (5'h1a == io_rdAddr[4:0]) begin // @[RegFile.scala 27:19]
        rf__26 <= io_rdData; // @[RegFile.scala 27:19]
      end
    end
    if (reset) begin // @[RegFile.scala 24:19]
      rf__27 <= 64'h0; // @[RegFile.scala 24:19]
    end else if (io_rdEn & io_rdAddr != 32'h0) begin // @[RegFile.scala 26:41]
      if (5'h1b == io_rdAddr[4:0]) begin // @[RegFile.scala 27:19]
        rf__27 <= io_rdData; // @[RegFile.scala 27:19]
      end
    end
    if (reset) begin // @[RegFile.scala 24:19]
      rf__28 <= 64'h0; // @[RegFile.scala 24:19]
    end else if (io_rdEn & io_rdAddr != 32'h0) begin // @[RegFile.scala 26:41]
      if (5'h1c == io_rdAddr[4:0]) begin // @[RegFile.scala 27:19]
        rf__28 <= io_rdData; // @[RegFile.scala 27:19]
      end
    end
    if (reset) begin // @[RegFile.scala 24:19]
      rf__29 <= 64'h0; // @[RegFile.scala 24:19]
    end else if (io_rdEn & io_rdAddr != 32'h0) begin // @[RegFile.scala 26:41]
      if (5'h1d == io_rdAddr[4:0]) begin // @[RegFile.scala 27:19]
        rf__29 <= io_rdData; // @[RegFile.scala 27:19]
      end
    end
    if (reset) begin // @[RegFile.scala 24:19]
      rf__30 <= 64'h0; // @[RegFile.scala 24:19]
    end else if (io_rdEn & io_rdAddr != 32'h0) begin // @[RegFile.scala 26:41]
      if (5'h1e == io_rdAddr[4:0]) begin // @[RegFile.scala 27:19]
        rf__30 <= io_rdData; // @[RegFile.scala 27:19]
      end
    end
    if (reset) begin // @[RegFile.scala 24:19]
      rf__31 <= 64'h0; // @[RegFile.scala 24:19]
    end else if (io_rdEn & io_rdAddr != 32'h0) begin // @[RegFile.scala 26:41]
      if (5'h1f == io_rdAddr[4:0]) begin // @[RegFile.scala 27:19]
        rf__31 <= io_rdData; // @[RegFile.scala 27:19]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  rf__0 = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  rf__1 = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  rf__2 = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  rf__3 = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  rf__4 = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  rf__5 = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  rf__6 = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  rf__7 = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  rf__8 = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  rf__9 = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  rf__10 = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  rf__11 = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  rf__12 = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  rf__13 = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  rf__14 = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  rf__15 = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  rf__16 = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  rf__17 = _RAND_17[63:0];
  _RAND_18 = {2{`RANDOM}};
  rf__18 = _RAND_18[63:0];
  _RAND_19 = {2{`RANDOM}};
  rf__19 = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  rf__20 = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  rf__21 = _RAND_21[63:0];
  _RAND_22 = {2{`RANDOM}};
  rf__22 = _RAND_22[63:0];
  _RAND_23 = {2{`RANDOM}};
  rf__23 = _RAND_23[63:0];
  _RAND_24 = {2{`RANDOM}};
  rf__24 = _RAND_24[63:0];
  _RAND_25 = {2{`RANDOM}};
  rf__25 = _RAND_25[63:0];
  _RAND_26 = {2{`RANDOM}};
  rf__26 = _RAND_26[63:0];
  _RAND_27 = {2{`RANDOM}};
  rf__27 = _RAND_27[63:0];
  _RAND_28 = {2{`RANDOM}};
  rf__28 = _RAND_28[63:0];
  _RAND_29 = {2{`RANDOM}};
  rf__29 = _RAND_29[63:0];
  _RAND_30 = {2{`RANDOM}};
  rf__30 = _RAND_30[63:0];
  _RAND_31 = {2{`RANDOM}};
  rf__31 = _RAND_31[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ContrGen(
  input  [31:0] io_inst,
  output [2:0]  io_branch,
  output [2:0]  io_immOp,
  output        io_rdEn,
  output [4:0]  io_rdAddr,
  output        io_typeL,
  output [3:0]  io_csrOp,
  output        io_aluCtr_aluA,
  output [1:0]  io_aluCtr_aluB,
  output [3:0]  io_aluCtr_aluOp,
  output [1:0]  io_memCtr_memtoReg,
  output        io_memCtr_memWr,
  output [2:0]  io_memCtr_memOP,
  output        io_regCtrl_rs1En,
  output        io_regCtrl_rs2En,
  output [4:0]  io_regCtrl_rs1Addr,
  output [4:0]  io_regCtrl_rs2Addr
);
  wire [31:0] _instLui_T = io_inst & 32'h7f; // @[ContrGen.scala 26:26]
  wire  instLui = 32'h37 == _instLui_T; // @[ContrGen.scala 26:26]
  wire  instAuipc = 32'h17 == _instLui_T; // @[ContrGen.scala 27:26]
  wire  typeU = instLui | instAuipc; // @[ContrGen.scala 28:29]
  wire [31:0] _instAddi_T = io_inst & 32'h707f; // @[ContrGen.scala 31:26]
  wire  instAddi = 32'h13 == _instAddi_T; // @[ContrGen.scala 31:26]
  wire  instAndi = 32'h7013 == _instAddi_T; // @[ContrGen.scala 32:26]
  wire  instXori = 32'h4013 == _instAddi_T; // @[ContrGen.scala 33:26]
  wire  instOri = 32'h6013 == _instAddi_T; // @[ContrGen.scala 34:26]
  wire [31:0] _instSlli_T = io_inst & 32'hfc00707f; // @[ContrGen.scala 35:26]
  wire  instSlli = 32'h1013 == _instSlli_T; // @[ContrGen.scala 35:26]
  wire  instSrli = 32'h5013 == _instSlli_T; // @[ContrGen.scala 36:26]
  wire  instSrai = 32'h40005013 == _instSlli_T; // @[ContrGen.scala 37:26]
  wire  instSlti = 32'h2013 == _instAddi_T; // @[ContrGen.scala 38:26]
  wire  instSltiu = 32'h3013 == _instAddi_T; // @[ContrGen.scala 39:26]
  wire  instAddiw = 32'h1b == _instAddi_T; // @[ContrGen.scala 40:26]
  wire [31:0] _instSlliw_T = io_inst & 32'hfe00707f; // @[ContrGen.scala 41:26]
  wire  instSlliw = 32'h101b == _instSlliw_T; // @[ContrGen.scala 41:26]
  wire  instSrliw = 32'h501b == _instSlliw_T; // @[ContrGen.scala 42:26]
  wire  instSraiw = 32'h4000501b == _instSlliw_T; // @[ContrGen.scala 43:26]
  wire  instJalr = 32'h67 == _instAddi_T; // @[ContrGen.scala 44:26]
  wire  instLb = 32'h3 == _instAddi_T; // @[ContrGen.scala 45:26]
  wire  instLh = 32'h1003 == _instAddi_T; // @[ContrGen.scala 46:26]
  wire  instLw = 32'h2003 == _instAddi_T; // @[ContrGen.scala 47:26]
  wire  instLd = 32'h3003 == _instAddi_T; // @[ContrGen.scala 48:26]
  wire  instLbu = 32'h4003 == _instAddi_T; // @[ContrGen.scala 49:26]
  wire  instLhu = 32'h5003 == _instAddi_T; // @[ContrGen.scala 50:26]
  wire  instLwu = 32'h6003 == _instAddi_T; // @[ContrGen.scala 51:26]
  wire  csrrw = 32'h1073 == _instAddi_T; // @[ContrGen.scala 54:22]
  wire  csrrs = 32'h2073 == _instAddi_T; // @[ContrGen.scala 55:22]
  wire  csrrc = 32'h3073 == _instAddi_T; // @[ContrGen.scala 56:22]
  wire  csrrwi = 32'h5073 == _instAddi_T; // @[ContrGen.scala 57:22]
  wire  csrrsi = 32'h6073 == _instAddi_T; // @[ContrGen.scala 58:22]
  wire  csrrci = 32'h7073 == _instAddi_T; // @[ContrGen.scala 59:22]
  wire  ecall = 32'h73 == io_inst; // @[ContrGen.scala 61:22]
  wire  mret = 32'h30200073 == io_inst; // @[ContrGen.scala 62:22]
  wire  _typeL_T_1 = instLb | instLh | instLw; // @[ContrGen.scala 69:32]
  wire  _typeL_T_4 = instLb | instLh | instLw | instLd | instLbu | instLhu; // @[ContrGen.scala 69:63]
  wire  instJal = 32'h6f == _instLui_T; // @[ContrGen.scala 73:26]
  wire  typeJ = instJal | instJalr; // @[ContrGen.scala 74:29]
  wire  instAdd = 32'h33 == _instSlliw_T; // @[ContrGen.scala 77:26]
  wire  instSub = 32'h40000033 == _instSlliw_T; // @[ContrGen.scala 78:26]
  wire  instSll = 32'h1033 == _instSlliw_T; // @[ContrGen.scala 79:26]
  wire  instSlt = 32'h2033 == _instSlliw_T; // @[ContrGen.scala 80:26]
  wire  instSltu = 32'h3033 == _instSlliw_T; // @[ContrGen.scala 81:26]
  wire  instXor = 32'h4033 == _instSlliw_T; // @[ContrGen.scala 82:26]
  wire  instSrl = 32'h5033 == _instSlliw_T; // @[ContrGen.scala 83:26]
  wire  instSra = 32'h40005033 == _instSlliw_T; // @[ContrGen.scala 84:26]
  wire  instOr = 32'h6033 == _instSlliw_T; // @[ContrGen.scala 85:26]
  wire  instAnd = 32'h7033 == _instSlliw_T; // @[ContrGen.scala 86:26]
  wire  instAddw = 32'h3b == _instSlliw_T; // @[ContrGen.scala 87:26]
  wire  instSubw = 32'h4000003b == _instSlliw_T; // @[ContrGen.scala 88:26]
  wire  instSllw = 32'h103b == _instSlliw_T; // @[ContrGen.scala 89:26]
  wire  instSrlw = 32'h503b == _instSlliw_T; // @[ContrGen.scala 90:26]
  wire  instSraw = 32'h4000503b == _instSlliw_T; // @[ContrGen.scala 91:26]
  wire  aluRem = 32'h200603b == _instSlliw_T; // @[ContrGen.scala 92:26]
  wire  instDiv = 32'h2004033 == _instSlliw_T; // @[ContrGen.scala 93:26]
  wire  instDivw = 32'h200403b == _instSlliw_T; // @[ContrGen.scala 94:26]
  wire  instMul = 32'h2000033 == _instSlliw_T; // @[ContrGen.scala 95:26]
  wire  instMulw = 32'h200003b == _instSlliw_T; // @[ContrGen.scala 96:26]
  wire  _typeR_T_4 = instAdd | instSub | instSll | instSlt | instSltu | instXor; // @[ContrGen.scala 97:78]
  wire  _typeR_T_9 = _typeR_T_4 | instSrl | instSra | instOr | instAnd | instAddw; // @[ContrGen.scala 98:78]
  wire  _typeR_T_14 = _typeR_T_9 | instSubw | instSllw | instSrlw | instSraw | aluRem; // @[ContrGen.scala 99:78]
  wire  typeR = _typeR_T_14 | instDiv | instDivw | instMul | instMulw | mret; // @[ContrGen.scala 100:78]
  wire  instBeq = 32'h63 == _instAddi_T; // @[ContrGen.scala 104:27]
  wire  instBne = 32'h1063 == _instAddi_T; // @[ContrGen.scala 105:27]
  wire  instBlt = 32'h4063 == _instAddi_T; // @[ContrGen.scala 106:27]
  wire  instBge = 32'h5063 == _instAddi_T; // @[ContrGen.scala 107:27]
  wire  instBltu = 32'h6063 == _instAddi_T; // @[ContrGen.scala 108:27]
  wire  instBgeu = 32'h7063 == _instAddi_T; // @[ContrGen.scala 109:27]
  wire  _typeB_T = instBeq | instBne; // @[ContrGen.scala 110:30]
  wire  typeB = instBeq | instBne | instBlt | instBge | instBltu | instBgeu; // @[ContrGen.scala 110:74]
  wire  instSb = 32'h23 == _instAddi_T; // @[ContrGen.scala 113:27]
  wire  instSh = 32'h1023 == _instAddi_T; // @[ContrGen.scala 114:27]
  wire  instSw = 32'h2023 == _instAddi_T; // @[ContrGen.scala 115:27]
  wire  instSd = 32'h3023 == _instAddi_T; // @[ContrGen.scala 116:27]
  wire  _typeS_T_1 = instSb | instSh | instSw; // @[ContrGen.scala 117:39]
  wire  typeS = instSb | instSh | instSw | instSd; // @[ContrGen.scala 117:49]
  wire  Ebreak = 32'h100073 == io_inst; // @[ContrGen.scala 120:21]
  wire  my_inst = 32'h7b == io_inst; // @[ContrGen.scala 123:22]
  wire  _typeW_T_3 = instAddw | instSubw | instSllw | instSlliw | instSraw; // @[ContrGen.scala 126:68]
  wire  _typeW_T_9 = _typeW_T_3 | instSrlw | instSrliw | instSraiw | instAddiw | aluRem | instDivw; // @[ContrGen.scala 127:76]
  wire  typeW = _typeW_T_9 | instMulw; // @[ContrGen.scala 128:14]
  wire  _io_aluCtr_aluB_T = typeR | typeB; // @[ContrGen.scala 134:12]
  wire [1:0] _io_aluCtr_aluB_T_1 = typeJ ? 2'h2 : 2'h1; // @[Mux.scala 101:16]
  wire  aluSub = instSub | instSubw; // @[ContrGen.scala 141:28]
  wire  aluSlt = instSlti | instSlt; // @[ContrGen.scala 142:29]
  wire  aluSltu = instSltiu | instSltu; // @[ContrGen.scala 143:29]
  wire  aluAnd = instAndi | instAnd; // @[ContrGen.scala 144:29]
  wire  aluOr = instOri | instOr; // @[ContrGen.scala 145:29]
  wire  aluXor = instXori | instXor; // @[ContrGen.scala 146:29]
  wire  aluSll = instSlli | instSlliw | instSll | instSllw; // @[ContrGen.scala 147:53]
  wire  aluSrl = instSrli | instSrliw | instSrl | instSrlw; // @[ContrGen.scala 148:53]
  wire  aluSra = instSrai | instSraiw | instSra | instSraw; // @[ContrGen.scala 149:53]
  wire  aluDiv = instDiv | instDivw; // @[ContrGen.scala 151:27]
  wire  aluMul = instMul | instMulw; // @[ContrGen.scala 152:27]
  wire  _io_aluCtr_aluOp_T_2 = aluSlt | instBlt | instBge; // @[ContrGen.scala 158:37]
  wire  _io_aluCtr_aluOp_T_6 = aluSltu | instBltu | instBgeu; // @[ContrGen.scala 160:40]
  wire [2:0] _io_aluCtr_aluOp_T_7 = aluAnd ? 3'h7 : 3'h0; // @[Mux.scala 101:16]
  wire [3:0] _io_aluCtr_aluOp_T_8 = aluMul ? 4'he : {{1'd0}, _io_aluCtr_aluOp_T_7}; // @[Mux.scala 101:16]
  wire [3:0] _io_aluCtr_aluOp_T_9 = aluOr ? 4'h6 : _io_aluCtr_aluOp_T_8; // @[Mux.scala 101:16]
  wire [3:0] _io_aluCtr_aluOp_T_10 = aluSra ? 4'hd : _io_aluCtr_aluOp_T_9; // @[Mux.scala 101:16]
  wire [3:0] _io_aluCtr_aluOp_T_11 = aluSrl ? 4'h5 : _io_aluCtr_aluOp_T_10; // @[Mux.scala 101:16]
  wire [3:0] _io_aluCtr_aluOp_T_12 = aluDiv ? 4'hc : _io_aluCtr_aluOp_T_11; // @[Mux.scala 101:16]
  wire [3:0] _io_aluCtr_aluOp_T_13 = aluXor ? 4'h4 : _io_aluCtr_aluOp_T_12; // @[Mux.scala 101:16]
  wire [3:0] _io_aluCtr_aluOp_T_14 = aluRem ? 4'hb : _io_aluCtr_aluOp_T_13; // @[Mux.scala 101:16]
  wire [3:0] _io_aluCtr_aluOp_T_15 = instLui ? 4'h3 : _io_aluCtr_aluOp_T_14; // @[Mux.scala 101:16]
  wire [3:0] _io_aluCtr_aluOp_T_16 = _io_aluCtr_aluOp_T_6 ? 4'ha : _io_aluCtr_aluOp_T_15; // @[Mux.scala 101:16]
  wire [3:0] _io_aluCtr_aluOp_T_17 = _typeB_T ? 4'h9 : _io_aluCtr_aluOp_T_16; // @[Mux.scala 101:16]
  wire [3:0] _io_aluCtr_aluOp_T_18 = _io_aluCtr_aluOp_T_2 ? 4'h2 : _io_aluCtr_aluOp_T_17; // @[Mux.scala 101:16]
  wire [3:0] _io_aluCtr_aluOp_T_19 = aluSll ? 4'h1 : _io_aluCtr_aluOp_T_18; // @[Mux.scala 101:16]
  wire  _io_branch_T = instBlt | instBltu; // @[ContrGen.scala 177:20]
  wire  _io_branch_T_1 = instBge | instBgeu; // @[ContrGen.scala 178:20]
  wire [2:0] _io_branch_T_2 = _io_branch_T_1 ? 3'h7 : 3'h0; // @[Mux.scala 101:16]
  wire [2:0] _io_branch_T_3 = _io_branch_T ? 3'h6 : _io_branch_T_2; // @[Mux.scala 101:16]
  wire [2:0] _io_branch_T_4 = instBne ? 3'h5 : _io_branch_T_3; // @[Mux.scala 101:16]
  wire [2:0] _io_branch_T_5 = instBeq ? 3'h4 : _io_branch_T_4; // @[Mux.scala 101:16]
  wire [2:0] _io_branch_T_6 = ecall ? 3'h3 : _io_branch_T_5; // @[Mux.scala 101:16]
  wire [2:0] _io_branch_T_7 = instJalr ? 3'h2 : _io_branch_T_6; // @[Mux.scala 101:16]
  wire  wRegEn = ~(typeS | typeB | Ebreak); // @[ContrGen.scala 185:16]
  wire  _io_immOp_T_8 = instAddi | instAddiw | instSlti | instSltiu | instXori | instOri | instAndi | instSlli |
    instSlliw | instSrli; // @[ContrGen.scala 190:120]
  wire  _io_immOp_T_15 = _io_immOp_T_8 | instSrliw | instSrai | instSraiw | instJalr | instLb | instLh | instLw; // @[ContrGen.scala 191:92]
  wire  _io_immOp_T_19 = _io_immOp_T_15 | instLwu | instLd | instLbu | instLhu; // @[ContrGen.scala 192:57]
  wire  _io_immOp_T_20 = instAuipc | instLui; // @[ContrGen.scala 193:22]
  wire  _io_immOp_T_23 = instSd | instSb | instSw | instSh; // @[ContrGen.scala 194:39]
  wire [2:0] _io_immOp_T_29 = instJal ? 3'h4 : 3'h7; // @[Mux.scala 101:16]
  wire [2:0] _io_immOp_T_30 = typeB ? 3'h3 : _io_immOp_T_29; // @[Mux.scala 101:16]
  wire [2:0] _io_immOp_T_31 = _io_immOp_T_23 ? 3'h2 : _io_immOp_T_30; // @[Mux.scala 101:16]
  wire [2:0] _io_immOp_T_32 = _io_immOp_T_20 ? 3'h1 : _io_immOp_T_31; // @[Mux.scala 101:16]
  wire  _io_memCtr_memtoReg_T_5 = _typeL_T_1 | instLwu | instLd | instLbu | instLhu; // @[ContrGen.scala 199:65]
  wire [1:0] _io_memCtr_memtoReg_T_6 = typeW ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire  _io_memCtr_memOP_T = instLb | instSb; // @[ContrGen.scala 205:19]
  wire  _io_memCtr_memOP_T_1 = instLh | instSh; // @[ContrGen.scala 206:19]
  wire  _io_memCtr_memOP_T_2 = instLw | instSw; // @[ContrGen.scala 207:19]
  wire  _io_memCtr_memOP_T_3 = instLd | instSd; // @[ContrGen.scala 208:19]
  wire [2:0] _io_memCtr_memOP_T_4 = instLwu ? 3'h6 : 3'h7; // @[Mux.scala 101:16]
  wire [2:0] _io_memCtr_memOP_T_5 = instLhu ? 3'h5 : _io_memCtr_memOP_T_4; // @[Mux.scala 101:16]
  wire [2:0] _io_memCtr_memOP_T_6 = instLbu ? 3'h4 : _io_memCtr_memOP_T_5; // @[Mux.scala 101:16]
  wire [2:0] _io_memCtr_memOP_T_7 = _io_memCtr_memOP_T_3 ? 3'h3 : _io_memCtr_memOP_T_6; // @[Mux.scala 101:16]
  wire [2:0] _io_memCtr_memOP_T_8 = _io_memCtr_memOP_T_2 ? 3'h2 : _io_memCtr_memOP_T_7; // @[Mux.scala 101:16]
  wire [2:0] _io_memCtr_memOP_T_9 = _io_memCtr_memOP_T_1 ? 3'h1 : _io_memCtr_memOP_T_8; // @[Mux.scala 101:16]
  wire [3:0] _io_csrOp_T = mret ? 4'h9 : 4'h0; // @[Mux.scala 101:16]
  wire [3:0] _io_csrOp_T_1 = ecall ? 4'h8 : _io_csrOp_T; // @[Mux.scala 101:16]
  wire [3:0] _io_csrOp_T_2 = csrrci ? 4'h7 : _io_csrOp_T_1; // @[Mux.scala 101:16]
  wire [3:0] _io_csrOp_T_3 = csrrsi ? 4'h6 : _io_csrOp_T_2; // @[Mux.scala 101:16]
  wire [3:0] _io_csrOp_T_4 = csrrwi ? 4'h5 : _io_csrOp_T_3; // @[Mux.scala 101:16]
  wire [3:0] _io_csrOp_T_5 = csrrc ? 4'h3 : _io_csrOp_T_4; // @[Mux.scala 101:16]
  wire [3:0] _io_csrOp_T_6 = csrrs ? 4'h2 : _io_csrOp_T_5; // @[Mux.scala 101:16]
  assign io_branch = instJal ? 3'h1 : _io_branch_T_7; // @[Mux.scala 101:16]
  assign io_immOp = _io_immOp_T_19 ? 3'h0 : _io_immOp_T_32; // @[Mux.scala 101:16]
  assign io_rdEn = ~(typeS | typeB | Ebreak); // @[ContrGen.scala 185:16]
  assign io_rdAddr = wRegEn ? io_inst[11:7] : 5'h0; // @[ContrGen.scala 187:19]
  assign io_typeL = _typeL_T_4 | instLwu; // @[ContrGen.scala 70:22]
  assign io_csrOp = csrrw ? 4'h1 : _io_csrOp_T_6; // @[Mux.scala 101:16]
  assign io_aluCtr_aluA = instAuipc | typeJ; // @[ContrGen.scala 131:35]
  assign io_aluCtr_aluB = _io_aluCtr_aluB_T ? 2'h0 : _io_aluCtr_aluB_T_1; // @[Mux.scala 101:16]
  assign io_aluCtr_aluOp = aluSub ? 4'h8 : _io_aluCtr_aluOp_T_19; // @[Mux.scala 101:16]
  assign io_memCtr_memtoReg = _io_memCtr_memtoReg_T_5 ? 2'h1 : _io_memCtr_memtoReg_T_6; // @[Mux.scala 101:16]
  assign io_memCtr_memWr = _typeS_T_1 | instSd; // @[ContrGen.scala 203:56]
  assign io_memCtr_memOP = _io_memCtr_memOP_T ? 3'h0 : _io_memCtr_memOP_T_9; // @[Mux.scala 101:16]
  assign io_regCtrl_rs1En = ~(typeU | instJal); // @[ContrGen.scala 180:23]
  assign io_regCtrl_rs2En = _io_aluCtr_aluB_T | typeS; // @[ContrGen.scala 181:40]
  assign io_regCtrl_rs1Addr = Ebreak | my_inst ? 5'ha : io_inst[19:15]; // @[ContrGen.scala 182:28]
  assign io_regCtrl_rs2Addr = io_inst[24:20]; // @[ContrGen.scala 183:29]
endmodule
module Decode(
  input         clock,
  input         reset,
  input         io_rdEn,
  input  [4:0]  io_rdAddr,
  input  [63:0] io_rdData,
  input         io_preRs1En,
  input  [4:0]  io_preRs1Addr,
  output [63:0] io_preRs1Data,
  output [63:0] io_preRs1x1Data,
  input         io_in_valid,
  input  [31:0] io_in_pc,
  input  [31:0] io_in_inst,
  input         io_in_takenPre,
  input  [31:0] io_in_takenPrePC,
  input         io_exeRdEn,
  input  [4:0]  io_exeRdAddr,
  input  [63:0] io_exeRdData,
  input         io_memRdEn,
  input  [4:0]  io_memRdAddr,
  input  [63:0] io_memRdData,
  input         io_wbRdEn,
  input  [4:0]  io_wbRdAddr,
  input  [63:0] io_wbRdData,
  output        io_bubbleId,
  output        io_sBubbleEx,
  output        io_sBubbleMem,
  output        io_out_valid,
  output [31:0] io_out_pc,
  output [31:0] io_out_inst,
  output        io_out_typeL,
  output        io_out_aluA,
  output [1:0]  io_out_aluB,
  output [3:0]  io_out_aluOp,
  output [2:0]  io_out_branch,
  output [1:0]  io_out_memtoReg,
  output        io_out_memWr,
  output [2:0]  io_out_memOp,
  output        io_out_rdEn,
  output [4:0]  io_out_rdAddr,
  output [63:0] io_out_rs1Data,
  output [63:0] io_out_rs2Data,
  output [63:0] io_out_imm,
  output [3:0]  io_out_csrOp,
  output        io_out_takenPre,
  output [31:0] io_out_takenPrePC,
  output [63:0] rf_10
);
  wire  regs_clock; // @[Decode.scala 43:20]
  wire  regs_reset; // @[Decode.scala 43:20]
  wire [63:0] regs_io_rs1Data; // @[Decode.scala 43:20]
  wire [63:0] regs_io_rs2Data; // @[Decode.scala 43:20]
  wire  regs_io_rdEn; // @[Decode.scala 43:20]
  wire [31:0] regs_io_rdAddr; // @[Decode.scala 43:20]
  wire [63:0] regs_io_rdData; // @[Decode.scala 43:20]
  wire  regs_io_preRs1En; // @[Decode.scala 43:20]
  wire [4:0] regs_io_preRs1Addr; // @[Decode.scala 43:20]
  wire [63:0] regs_io_preRs1Data; // @[Decode.scala 43:20]
  wire [63:0] regs_io_preRs1x1Data; // @[Decode.scala 43:20]
  wire  regs_io_ctrl_rs1En; // @[Decode.scala 43:20]
  wire  regs_io_ctrl_rs2En; // @[Decode.scala 43:20]
  wire [4:0] regs_io_ctrl_rs1Addr; // @[Decode.scala 43:20]
  wire [4:0] regs_io_ctrl_rs2Addr; // @[Decode.scala 43:20]
  wire [63:0] regs_rf_10; // @[Decode.scala 43:20]
  wire [31:0] imm_io_inst; // @[Decode.scala 44:20]
  wire [2:0] imm_io_immOp; // @[Decode.scala 44:20]
  wire [63:0] imm_io_imm; // @[Decode.scala 44:20]
  wire [31:0] con_io_inst; // @[Decode.scala 45:20]
  wire [2:0] con_io_branch; // @[Decode.scala 45:20]
  wire [2:0] con_io_immOp; // @[Decode.scala 45:20]
  wire  con_io_rdEn; // @[Decode.scala 45:20]
  wire [4:0] con_io_rdAddr; // @[Decode.scala 45:20]
  wire  con_io_typeL; // @[Decode.scala 45:20]
  wire [3:0] con_io_csrOp; // @[Decode.scala 45:20]
  wire  con_io_aluCtr_aluA; // @[Decode.scala 45:20]
  wire [1:0] con_io_aluCtr_aluB; // @[Decode.scala 45:20]
  wire [3:0] con_io_aluCtr_aluOp; // @[Decode.scala 45:20]
  wire [1:0] con_io_memCtr_memtoReg; // @[Decode.scala 45:20]
  wire  con_io_memCtr_memWr; // @[Decode.scala 45:20]
  wire [2:0] con_io_memCtr_memOP; // @[Decode.scala 45:20]
  wire  con_io_regCtrl_rs1En; // @[Decode.scala 45:20]
  wire  con_io_regCtrl_rs2En; // @[Decode.scala 45:20]
  wire [4:0] con_io_regCtrl_rs1Addr; // @[Decode.scala 45:20]
  wire [4:0] con_io_regCtrl_rs2Addr; // @[Decode.scala 45:20]
  wire [4:0] rs1Addr = con_io_regCtrl_rs1En ? con_io_regCtrl_rs1Addr : 5'h0; // @[Decode.scala 63:20]
  wire [4:0] rs2Addr = con_io_regCtrl_rs2En ? con_io_regCtrl_rs2Addr : 5'h0; // @[Decode.scala 64:20]
  wire  _rdRs1HitEx_T_2 = rs1Addr != 5'h0; // @[Decode.scala 65:73]
  wire  rdRs1HitEx = io_exeRdEn & rs1Addr == io_exeRdAddr & rs1Addr != 5'h0; // @[Decode.scala 65:61]
  wire  rdRs1HitMem = io_memRdEn & rs1Addr == io_memRdAddr & _rdRs1HitEx_T_2; // @[Decode.scala 66:62]
  wire  rdRs1HitWb = io_wbRdEn & rs1Addr == io_wbRdAddr & _rdRs1HitEx_T_2; // @[Decode.scala 67:59]
  wire  _rdRs2HitEx_T_2 = rs2Addr != 5'h0; // @[Decode.scala 69:73]
  wire  rdRs2HitEx = io_exeRdEn & rs2Addr == io_exeRdAddr & rs2Addr != 5'h0; // @[Decode.scala 69:61]
  wire  rdRs2HitMem = io_memRdEn & rs2Addr == io_memRdAddr & _rdRs2HitEx_T_2; // @[Decode.scala 70:62]
  wire  rdRs2HitWb = io_wbRdEn & rs2Addr == io_wbRdAddr & _rdRs2HitEx_T_2; // @[Decode.scala 71:59]
  wire [63:0] _rs1Data_T = rdRs1HitWb ? io_wbRdData : regs_io_rs1Data; // @[Decode.scala 76:8]
  wire [63:0] _rs1Data_T_1 = rdRs1HitMem ? io_memRdData : _rs1Data_T; // @[Decode.scala 75:8]
  wire [63:0] _rs1Data_T_2 = rdRs1HitEx ? io_exeRdData : _rs1Data_T_1; // @[Decode.scala 74:8]
  wire [63:0] _rs2Data_T = rdRs2HitWb ? io_wbRdData : regs_io_rs2Data; // @[Decode.scala 81:8]
  wire [63:0] _rs2Data_T_1 = rdRs2HitMem ? io_memRdData : _rs2Data_T; // @[Decode.scala 80:8]
  wire [63:0] _rs2Data_T_2 = rdRs2HitEx ? io_exeRdData : _rs2Data_T_1; // @[Decode.scala 79:8]
  RegFile regs ( // @[Decode.scala 43:20]
    .clock(regs_clock),
    .reset(regs_reset),
    .io_rs1Data(regs_io_rs1Data),
    .io_rs2Data(regs_io_rs2Data),
    .io_rdEn(regs_io_rdEn),
    .io_rdAddr(regs_io_rdAddr),
    .io_rdData(regs_io_rdData),
    .io_preRs1En(regs_io_preRs1En),
    .io_preRs1Addr(regs_io_preRs1Addr),
    .io_preRs1Data(regs_io_preRs1Data),
    .io_preRs1x1Data(regs_io_preRs1x1Data),
    .io_ctrl_rs1En(regs_io_ctrl_rs1En),
    .io_ctrl_rs2En(regs_io_ctrl_rs2En),
    .io_ctrl_rs1Addr(regs_io_ctrl_rs1Addr),
    .io_ctrl_rs2Addr(regs_io_ctrl_rs2Addr),
    .rf_10(regs_rf_10)
  );
  ImmGen imm ( // @[Decode.scala 44:20]
    .io_inst(imm_io_inst),
    .io_immOp(imm_io_immOp),
    .io_imm(imm_io_imm)
  );
  ContrGen con ( // @[Decode.scala 45:20]
    .io_inst(con_io_inst),
    .io_branch(con_io_branch),
    .io_immOp(con_io_immOp),
    .io_rdEn(con_io_rdEn),
    .io_rdAddr(con_io_rdAddr),
    .io_typeL(con_io_typeL),
    .io_csrOp(con_io_csrOp),
    .io_aluCtr_aluA(con_io_aluCtr_aluA),
    .io_aluCtr_aluB(con_io_aluCtr_aluB),
    .io_aluCtr_aluOp(con_io_aluCtr_aluOp),
    .io_memCtr_memtoReg(con_io_memCtr_memtoReg),
    .io_memCtr_memWr(con_io_memCtr_memWr),
    .io_memCtr_memOP(con_io_memCtr_memOP),
    .io_regCtrl_rs1En(con_io_regCtrl_rs1En),
    .io_regCtrl_rs2En(con_io_regCtrl_rs2En),
    .io_regCtrl_rs1Addr(con_io_regCtrl_rs1Addr),
    .io_regCtrl_rs2Addr(con_io_regCtrl_rs2Addr)
  );
  assign io_preRs1Data = regs_io_preRs1Data; // @[Decode.scala 53:17]
  assign io_preRs1x1Data = regs_io_preRs1x1Data; // @[Decode.scala 54:19]
  assign io_bubbleId = rdRs1HitEx | rdRs2HitEx; // @[Decode.scala 129:30]
  assign io_sBubbleEx = rdRs1HitEx | rdRs2HitEx; // @[Decode.scala 132:31]
  assign io_sBubbleMem = rdRs1HitMem | rdRs2HitMem; // @[Decode.scala 133:33]
  assign io_out_valid = io_in_valid; // @[Decode.scala 104:19]
  assign io_out_pc = io_in_pc; // @[Decode.scala 105:19]
  assign io_out_inst = io_in_inst; // @[Decode.scala 106:19]
  assign io_out_typeL = con_io_typeL; // @[Decode.scala 107:19]
  assign io_out_aluA = con_io_aluCtr_aluA; // @[Decode.scala 108:19]
  assign io_out_aluB = con_io_aluCtr_aluB; // @[Decode.scala 109:19]
  assign io_out_aluOp = con_io_aluCtr_aluOp; // @[Decode.scala 110:19]
  assign io_out_branch = con_io_branch; // @[Decode.scala 111:19]
  assign io_out_memtoReg = con_io_memCtr_memtoReg; // @[Decode.scala 112:19]
  assign io_out_memWr = con_io_memCtr_memWr; // @[Decode.scala 113:19]
  assign io_out_memOp = con_io_memCtr_memOP; // @[Decode.scala 114:19]
  assign io_out_rdEn = con_io_rdEn; // @[Decode.scala 116:19]
  assign io_out_rdAddr = con_io_rdAddr; // @[Decode.scala 117:19]
  assign io_out_rs1Data = con_io_regCtrl_rs1En ? _rs1Data_T_2 : 64'h0; // @[Decode.scala 73:20]
  assign io_out_rs2Data = con_io_regCtrl_rs2En ? _rs2Data_T_2 : 64'h0; // @[Decode.scala 78:20]
  assign io_out_imm = imm_io_imm; // @[Decode.scala 120:19]
  assign io_out_csrOp = con_io_csrOp; // @[Decode.scala 125:19]
  assign io_out_takenPre = io_in_takenPre; // @[Decode.scala 126:19]
  assign io_out_takenPrePC = io_in_takenPrePC; // @[Decode.scala 127:21]
  assign rf_10 = regs_rf_10;
  assign regs_clock = clock;
  assign regs_reset = reset;
  assign regs_io_rdEn = io_rdEn; // @[Decode.scala 48:16]
  assign regs_io_rdAddr = {{27'd0}, io_rdAddr}; // @[Decode.scala 49:18]
  assign regs_io_rdData = io_rdData; // @[Decode.scala 50:18]
  assign regs_io_preRs1En = io_preRs1En; // @[Decode.scala 51:20]
  assign regs_io_preRs1Addr = io_preRs1Addr; // @[Decode.scala 52:22]
  assign regs_io_ctrl_rs1En = con_io_regCtrl_rs1En; // @[Decode.scala 47:16]
  assign regs_io_ctrl_rs2En = con_io_regCtrl_rs2En; // @[Decode.scala 47:16]
  assign regs_io_ctrl_rs1Addr = con_io_regCtrl_rs1Addr; // @[Decode.scala 47:16]
  assign regs_io_ctrl_rs2Addr = con_io_regCtrl_rs2Addr; // @[Decode.scala 47:16]
  assign imm_io_inst = io_in_inst; // @[Decode.scala 56:15]
  assign imm_io_immOp = con_io_immOp; // @[Decode.scala 57:16]
  assign con_io_inst = io_in_inst; // @[Decode.scala 58:15]
endmodule
module ALU(
  input  [1:0]  io_memtoReg,
  input  [31:0] io_pc,
  output [63:0] io_aluRes,
  output        io_less,
  output        io_zero,
  input         ctrl_aluA,
  input  [1:0]  ctrl_aluB,
  input  [3:0]  ctrl_aluOp,
  input  [63:0] data_rData1,
  input  [63:0] data_rData2,
  input  [63:0] data_imm
);
  wire [63:0] Asrc = ~ctrl_aluA ? data_rData1 : {{32'd0}, io_pc}; // @[ALU.scala 23:19]
  wire  instW = io_memtoReg[1]; // @[ALU.scala 25:28]
  wire  in1_signBit = Asrc[31]; // @[BitUtils.scala 18:20]
  wire [31:0] _in1_T_3 = in1_signBit ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _in1_T_4 = {_in1_T_3,Asrc[31:0]}; // @[Cat.scala 31:58]
  wire [63:0] _in1_T_6 = {32'h0,Asrc[31:0]}; // @[Cat.scala 31:58]
  wire [63:0] _in1_T_7 = ctrl_aluOp == 4'hd ? _in1_T_4 : _in1_T_6; // @[ALU.scala 26:30]
  wire [63:0] in1 = instW ? _in1_T_7 : Asrc; // @[ALU.scala 26:18]
  wire [63:0] _in2_T_1 = 2'h1 == ctrl_aluB ? data_imm : data_rData2; // @[Mux.scala 81:58]
  wire [63:0] _in2_T_3 = 2'h2 == ctrl_aluB ? 64'h4 : _in2_T_1; // @[Mux.scala 81:58]
  wire [63:0] in2 = 2'h3 == ctrl_aluB ? 64'h0 : _in2_T_3; // @[Mux.scala 81:58]
  wire [5:0] shamt = instW ? {{1'd0}, in2[4:0]} : in2[5:0]; // @[ALU.scala 36:20]
  wire [63:0] addRes = in1 + in2; // @[ALU.scala 38:25]
  wire [63:0] subRes = in1 - in2; // @[ALU.scala 39:25]
  wire [63:0] xorRes = in1 ^ in2; // @[ALU.scala 40:25]
  wire [63:0] orRes = in1 | in2; // @[ALU.scala 41:25]
  wire [63:0] andRes = in1 & in2; // @[ALU.scala 42:25]
  wire [126:0] _GEN_0 = {{63'd0}, in1}; // @[ALU.scala 43:28]
  wire [126:0] _sLRes_T = _GEN_0 << shamt; // @[ALU.scala 43:28]
  wire [63:0] sLRes = _sLRes_T[63:0]; // @[ALU.scala 43:37]
  wire [63:0] sRLRes = in1 >> shamt; // @[ALU.scala 44:27]
  wire [63:0] _sRARes_T = instW ? _in1_T_7 : Asrc; // @[ALU.scala 45:33]
  wire [63:0] sRARes = $signed(_sRARes_T) >>> shamt; // @[ALU.scala 45:52]
  wire [63:0] _sLTRes_T_1 = 2'h3 == ctrl_aluB ? 64'h0 : _in2_T_3; // @[ALU.scala 47:48]
  wire  sLTRes = $signed(_sRARes_T) < $signed(_sLTRes_T_1); // @[ALU.scala 47:36]
  wire  sLTURes = in1 < in2; // @[ALU.scala 48:27]
  wire [63:0] remwRes = $signed(_sRARes_T) % $signed(_sLTRes_T_1); // @[ALU.scala 50:48]
  wire [63:0] divRes = in1 / in2; // @[ALU.scala 51:27]
  wire [127:0] mulRes = in1 * in2; // @[ALU.scala 52:27]
  wire [63:0] _aluResult_T_1 = 4'h0 == ctrl_aluOp ? addRes : 64'h0; // @[Mux.scala 81:58]
  wire [63:0] _aluResult_T_3 = 4'h8 == ctrl_aluOp ? subRes : _aluResult_T_1; // @[Mux.scala 81:58]
  wire [63:0] _aluResult_T_5 = 4'h9 == ctrl_aluOp ? subRes : _aluResult_T_3; // @[Mux.scala 81:58]
  wire [63:0] _aluResult_T_7 = 4'h2 == ctrl_aluOp ? {{63'd0}, sLTRes} : _aluResult_T_5; // @[Mux.scala 81:58]
  wire [63:0] _aluResult_T_9 = 4'ha == ctrl_aluOp ? {{63'd0}, sLTURes} : _aluResult_T_7; // @[Mux.scala 81:58]
  wire [63:0] _aluResult_T_11 = 4'h5 == ctrl_aluOp ? sRLRes : _aluResult_T_9; // @[Mux.scala 81:58]
  wire [63:0] _aluResult_T_13 = 4'hd == ctrl_aluOp ? sRARes : _aluResult_T_11; // @[Mux.scala 81:58]
  wire [63:0] _aluResult_T_15 = 4'h1 == ctrl_aluOp ? sLRes : _aluResult_T_13; // @[Mux.scala 81:58]
  wire [63:0] _aluResult_T_17 = 4'h3 == ctrl_aluOp ? in2 : _aluResult_T_15; // @[Mux.scala 81:58]
  wire [63:0] _aluResult_T_19 = 4'hb == ctrl_aluOp ? remwRes : _aluResult_T_17; // @[Mux.scala 81:58]
  wire [63:0] _aluResult_T_21 = 4'h4 == ctrl_aluOp ? xorRes : _aluResult_T_19; // @[Mux.scala 81:58]
  wire [63:0] _aluResult_T_23 = 4'hc == ctrl_aluOp ? divRes : _aluResult_T_21; // @[Mux.scala 81:58]
  wire [63:0] _aluResult_T_25 = 4'h6 == ctrl_aluOp ? orRes : _aluResult_T_23; // @[Mux.scala 81:58]
  wire [127:0] _aluResult_T_27 = 4'he == ctrl_aluOp ? mulRes : {{64'd0}, _aluResult_T_25}; // @[Mux.scala 81:58]
  wire [127:0] aluResult = 4'h7 == ctrl_aluOp ? {{64'd0}, andRes} : _aluResult_T_27; // @[Mux.scala 81:58]
  wire  io_aluRes_signBit = aluResult[31]; // @[BitUtils.scala 18:20]
  wire [31:0] _io_aluRes_T_2 = io_aluRes_signBit ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _io_aluRes_T_3 = {_io_aluRes_T_2,aluResult[31:0]}; // @[Cat.scala 31:58]
  wire [127:0] _io_aluRes_T_4 = instW ? {{64'd0}, _io_aluRes_T_3} : aluResult; // @[ALU.scala 80:21]
  assign io_aluRes = _io_aluRes_T_4[63:0]; // @[ALU.scala 80:15]
  assign io_less = ctrl_aluOp[3] ? sLTURes : sLTRes; // @[ALU.scala 78:19]
  assign io_zero = aluResult == 128'h0; // @[ALU.scala 79:27]
endmodule
module NextPC(
  input  [31:0] io_pc,
  input  [63:0] io_imm,
  input  [63:0] io_rs1Data,
  input  [2:0]  io_branch,
  input         io_less,
  input         io_zero,
  input         io_exc,
  input  [3:0]  io_csrOp,
  input  [63:0] io_mepc,
  input  [63:0] io_mtvec,
  input         io_time_int,
  output [31:0] io_nextPC,
  output [1:0]  io_pcSrc
);
  wire  less = io_branch == 3'h7 ? ~io_less : io_less; // @[NextPC.scala 29:17]
  wire [3:0] _pcSrc_T_1 = {io_branch,io_zero}; // @[NextPC.scala 32:43]
  wire [3:0] _pcSrc_T_7 = {io_branch,less}; // @[NextPC.scala 33:20]
  wire  _pcSrc_T_8 = _pcSrc_T_7 == 4'hc; // @[NextPC.scala 33:28]
  wire  _pcSrc_T_9 = io_branch == 3'h0 | _pcSrc_T_1 == 4'h8 | _pcSrc_T_1 == 4'hb | _pcSrc_T_8; // @[NextPC.scala 32:109]
  wire  _pcSrc_T_12 = _pcSrc_T_9 | _pcSrc_T_7 == 4'he; // @[NextPC.scala 33:43]
  wire  _pcSrc_T_21 = _pcSrc_T_7 == 4'hd; // @[NextPC.scala 35:28]
  wire  _pcSrc_T_22 = io_branch == 3'h1 | _pcSrc_T_1 == 4'h9 | _pcSrc_T_1 == 4'ha | _pcSrc_T_21; // @[NextPC.scala 34:108]
  wire  _pcSrc_T_25 = _pcSrc_T_22 | _pcSrc_T_7 == 4'hf; // @[NextPC.scala 35:43]
  wire  _pcSrc_T_28 = io_branch == 3'h2 | io_branch == 3'h3; // @[NextPC.scala 36:31]
  wire [1:0] _pcSrc_T_29 = _pcSrc_T_28 ? 2'h3 : 2'h1; // @[Mux.scala 101:16]
  wire [1:0] _pcSrc_T_30 = _pcSrc_T_25 ? 2'h2 : _pcSrc_T_29; // @[Mux.scala 101:16]
  wire [1:0] pcSrc = _pcSrc_T_12 ? 2'h0 : _pcSrc_T_30; // @[Mux.scala 101:16]
  wire [31:0] _GEN_0 = {io_mtvec[31:2], 2'h0}; // @[NextPC.scala 40:63]
  wire [32:0] _io_nextPC_T_4 = {{1'd0}, _GEN_0}; // @[NextPC.scala 40:63]
  wire [63:0] _io_nextPC_T_5 = ~io_csrOp[0] | io_time_int ? {{31'd0}, _io_nextPC_T_4} : io_mepc; // @[NextPC.scala 40:8]
  wire [31:0] _io_nextPC_T_7 = io_pc + 32'h4; // @[NextPC.scala 42:25]
  wire [63:0] _GEN_1 = {{32'd0}, io_pc}; // @[NextPC.scala 43:25]
  wire [63:0] _io_nextPC_T_9 = _GEN_1 + io_imm; // @[NextPC.scala 43:25]
  wire [63:0] _io_nextPC_T_11 = io_rs1Data + io_imm; // @[NextPC.scala 44:30]
  wire [31:0] _io_nextPC_T_13 = 2'h0 == pcSrc ? _io_nextPC_T_7 : 32'h80000000; // @[Mux.scala 81:58]
  wire [63:0] _io_nextPC_T_15 = 2'h2 == pcSrc ? _io_nextPC_T_9 : {{32'd0}, _io_nextPC_T_13}; // @[Mux.scala 81:58]
  wire [63:0] _io_nextPC_T_17 = 2'h3 == pcSrc ? _io_nextPC_T_11 : _io_nextPC_T_15; // @[Mux.scala 81:58]
  wire [63:0] _io_nextPC_T_18 = io_exc ? _io_nextPC_T_5 : _io_nextPC_T_17; // @[NextPC.scala 39:19]
  assign io_nextPC = _io_nextPC_T_18[31:0]; // @[NextPC.scala 39:13]
  assign io_pcSrc = _pcSrc_T_12 ? 2'h0 : _pcSrc_T_30; // @[Mux.scala 101:16]
endmodule
module Execution(
  input         io_in_valid,
  input  [31:0] io_in_pc,
  input  [31:0] io_in_inst,
  input         io_in_typeL,
  input         io_in_aluA,
  input  [1:0]  io_in_aluB,
  input  [3:0]  io_in_aluOp,
  input  [2:0]  io_in_branch,
  input  [1:0]  io_in_memtoReg,
  input         io_in_memWr,
  input  [2:0]  io_in_memOp,
  input         io_in_rdEn,
  input  [4:0]  io_in_rdAddr,
  input  [63:0] io_in_rs1Data,
  input  [63:0] io_in_rs2Data,
  input  [63:0] io_in_imm,
  input  [3:0]  io_in_csrOp,
  input         io_in_takenPre,
  input  [31:0] io_in_takenPrePC,
  output        io_out_valid,
  output [31:0] io_out_pc,
  output [31:0] io_out_inst,
  output        io_out_typeL,
  output        io_out_aluA,
  output [1:0]  io_out_aluB,
  output [3:0]  io_out_aluOp,
  output [2:0]  io_out_branch,
  output [1:0]  io_out_memtoReg,
  output        io_out_memWr,
  output [2:0]  io_out_memOp,
  output        io_out_rdEn,
  output [4:0]  io_out_rdAddr,
  output [63:0] io_out_rs1Data,
  output [63:0] io_out_rs2Data,
  output [63:0] io_out_imm,
  output [31:0] io_out_nextPC,
  output [63:0] io_out_aluRes,
  output [3:0]  io_out_csrOp,
  output        io_out_takenPre,
  output [31:0] io_out_takenPrePC,
  output [63:0] io_exeRdData,
  output        io_bubbleEx,
  output        io_takenValid,
  output        io_takenValidJalr,
  output        io_takenMiss,
  output        io_exTakenPre,
  output [31:0] io_takenPC,
  output        io_exeX1En,
  output [63:0] io_exeAluRes,
  input         io_exc,
  input  [3:0]  io_csrOp,
  input  [63:0] io_mepc,
  input  [63:0] io_mtvec,
  input         io_time_int
);
  wire [1:0] alu_io_memtoReg; // @[Execution.scala 27:21]
  wire [31:0] alu_io_pc; // @[Execution.scala 27:21]
  wire [63:0] alu_io_aluRes; // @[Execution.scala 27:21]
  wire  alu_io_less; // @[Execution.scala 27:21]
  wire  alu_io_zero; // @[Execution.scala 27:21]
  wire  alu_ctrl_aluA; // @[Execution.scala 27:21]
  wire [1:0] alu_ctrl_aluB; // @[Execution.scala 27:21]
  wire [3:0] alu_ctrl_aluOp; // @[Execution.scala 27:21]
  wire [63:0] alu_data_rData1; // @[Execution.scala 27:21]
  wire [63:0] alu_data_rData2; // @[Execution.scala 27:21]
  wire [63:0] alu_data_imm; // @[Execution.scala 27:21]
  wire [31:0] nextPC_io_pc; // @[Execution.scala 28:24]
  wire [63:0] nextPC_io_imm; // @[Execution.scala 28:24]
  wire [63:0] nextPC_io_rs1Data; // @[Execution.scala 28:24]
  wire [2:0] nextPC_io_branch; // @[Execution.scala 28:24]
  wire  nextPC_io_less; // @[Execution.scala 28:24]
  wire  nextPC_io_zero; // @[Execution.scala 28:24]
  wire  nextPC_io_exc; // @[Execution.scala 28:24]
  wire [3:0] nextPC_io_csrOp; // @[Execution.scala 28:24]
  wire [63:0] nextPC_io_mepc; // @[Execution.scala 28:24]
  wire [63:0] nextPC_io_mtvec; // @[Execution.scala 28:24]
  wire  nextPC_io_time_int; // @[Execution.scala 28:24]
  wire [31:0] nextPC_io_nextPC; // @[Execution.scala 28:24]
  wire [1:0] nextPC_io_pcSrc; // @[Execution.scala 28:24]
  ALU alu ( // @[Execution.scala 27:21]
    .io_memtoReg(alu_io_memtoReg),
    .io_pc(alu_io_pc),
    .io_aluRes(alu_io_aluRes),
    .io_less(alu_io_less),
    .io_zero(alu_io_zero),
    .ctrl_aluA(alu_ctrl_aluA),
    .ctrl_aluB(alu_ctrl_aluB),
    .ctrl_aluOp(alu_ctrl_aluOp),
    .data_rData1(alu_data_rData1),
    .data_rData2(alu_data_rData2),
    .data_imm(alu_data_imm)
  );
  NextPC nextPC ( // @[Execution.scala 28:24]
    .io_pc(nextPC_io_pc),
    .io_imm(nextPC_io_imm),
    .io_rs1Data(nextPC_io_rs1Data),
    .io_branch(nextPC_io_branch),
    .io_less(nextPC_io_less),
    .io_zero(nextPC_io_zero),
    .io_exc(nextPC_io_exc),
    .io_csrOp(nextPC_io_csrOp),
    .io_mepc(nextPC_io_mepc),
    .io_mtvec(nextPC_io_mtvec),
    .io_time_int(nextPC_io_time_int),
    .io_nextPC(nextPC_io_nextPC),
    .io_pcSrc(nextPC_io_pcSrc)
  );
  assign io_out_valid = io_in_valid; // @[Execution.scala 76:19]
  assign io_out_pc = io_in_pc; // @[Execution.scala 77:19]
  assign io_out_inst = io_in_inst; // @[Execution.scala 78:19]
  assign io_out_typeL = io_in_typeL; // @[Execution.scala 79:19]
  assign io_out_aluA = io_in_aluA; // @[Execution.scala 80:19]
  assign io_out_aluB = io_in_aluB; // @[Execution.scala 81:19]
  assign io_out_aluOp = io_in_aluOp; // @[Execution.scala 82:19]
  assign io_out_branch = io_in_branch; // @[Execution.scala 83:19]
  assign io_out_memtoReg = io_in_memtoReg; // @[Execution.scala 84:19]
  assign io_out_memWr = io_in_memWr; // @[Execution.scala 85:19]
  assign io_out_memOp = io_in_memOp; // @[Execution.scala 86:19]
  assign io_out_rdEn = io_in_rdEn; // @[Execution.scala 88:19]
  assign io_out_rdAddr = io_in_rdAddr; // @[Execution.scala 89:19]
  assign io_out_rs1Data = io_in_rs1Data; // @[Execution.scala 90:19]
  assign io_out_rs2Data = io_in_rs2Data; // @[Execution.scala 91:19]
  assign io_out_imm = io_in_imm; // @[Execution.scala 92:19]
  assign io_out_nextPC = nextPC_io_nextPC; // @[Execution.scala 94:19]
  assign io_out_aluRes = alu_io_aluRes; // @[Execution.scala 95:19]
  assign io_out_csrOp = io_in_csrOp; // @[Execution.scala 97:19]
  assign io_out_takenPre = io_in_takenPre; // @[Execution.scala 98:19]
  assign io_out_takenPrePC = io_in_takenPrePC; // @[Execution.scala 99:21]
  assign io_exeRdData = alu_io_aluRes; // @[Execution.scala 101:16]
  assign io_bubbleEx = io_in_typeL; // @[Execution.scala 102:15]
  assign io_takenValid = io_in_branch[2]; // @[Execution.scala 104:29]
  assign io_takenValidJalr = io_in_branch == 3'h2; // @[Execution.scala 105:35]
  assign io_takenMiss = io_in_takenPre ? io_in_takenPrePC != nextPC_io_nextPC : nextPC_io_pcSrc != 2'h0; // @[Execution.scala 106:23]
  assign io_exTakenPre = nextPC_io_pcSrc != 2'h0; // @[Execution.scala 107:29]
  assign io_takenPC = io_in_pc; // @[Execution.scala 108:17]
  assign io_exeX1En = io_in_rdEn & io_in_rdAddr == 5'h1; // @[Execution.scala 110:28]
  assign io_exeAluRes = alu_io_aluRes; // @[Execution.scala 111:16]
  assign alu_io_memtoReg = io_in_memtoReg; // @[Execution.scala 36:21]
  assign alu_io_pc = io_in_pc; // @[Execution.scala 37:15]
  assign alu_ctrl_aluA = io_in_aluA; // @[Execution.scala 30:25]
  assign alu_ctrl_aluB = io_in_aluB; // @[Execution.scala 31:25]
  assign alu_ctrl_aluOp = io_in_aluOp; // @[Execution.scala 32:26]
  assign alu_data_rData1 = io_in_rs1Data; // @[Execution.scala 33:27]
  assign alu_data_rData2 = io_in_rs2Data; // @[Execution.scala 34:27]
  assign alu_data_imm = io_in_imm; // @[Execution.scala 35:24]
  assign nextPC_io_pc = io_in_pc; // @[Execution.scala 39:18]
  assign nextPC_io_imm = io_in_imm; // @[Execution.scala 40:19]
  assign nextPC_io_rs1Data = io_in_rs1Data; // @[Execution.scala 41:23]
  assign nextPC_io_branch = io_in_branch; // @[Execution.scala 42:22]
  assign nextPC_io_less = alu_io_less; // @[Execution.scala 43:20]
  assign nextPC_io_zero = alu_io_zero; // @[Execution.scala 44:20]
  assign nextPC_io_exc = io_exc; // @[Execution.scala 46:19]
  assign nextPC_io_csrOp = io_csrOp; // @[Execution.scala 47:21]
  assign nextPC_io_mepc = io_mepc; // @[Execution.scala 48:20]
  assign nextPC_io_mtvec = io_mtvec; // @[Execution.scala 49:21]
  assign nextPC_io_time_int = io_time_int; // @[Execution.scala 50:24]
endmodule
module DataMem(
  input          clock,
  input          reset,
  output         io_dmem_data_valid,
  input          io_dmem_data_ready,
  output         io_dmem_data_req,
  output [31:0]  io_dmem_data_addr,
  output [1:0]   io_dmem_data_size,
  output [7:0]   io_dmem_data_strb,
  input  [63:0]  io_dmem_data_read,
  output [127:0] io_dmem_data_write,
  input          io_IFDone,
  input          io_in_valid,
  input  [31:0]  io_in_pc,
  input  [31:0]  io_in_inst,
  input          io_in_typeL,
  input          io_in_aluA,
  input  [1:0]   io_in_aluB,
  input  [3:0]   io_in_aluOp,
  input  [2:0]   io_in_branch,
  input  [1:0]   io_in_memtoReg,
  input          io_in_memWr,
  input  [2:0]   io_in_memOp,
  input          io_in_rdEn,
  input  [4:0]   io_in_rdAddr,
  input  [63:0]  io_in_rs1Data,
  input  [63:0]  io_in_rs2Data,
  input  [63:0]  io_in_imm,
  input  [63:0]  io_in_aluRes,
  input  [3:0]   io_in_csrOp,
  input          io_in_takenPre,
  input  [31:0]  io_in_takenPrePC,
  output         io_out_valid,
  output [31:0]  io_out_pc,
  output [31:0]  io_out_inst,
  output         io_out_typeL,
  output         io_out_aluA,
  output [1:0]   io_out_aluB,
  output [3:0]   io_out_aluOp,
  output [2:0]   io_out_branch,
  output [1:0]   io_out_memtoReg,
  output         io_out_memWr,
  output [2:0]   io_out_memOp,
  output [31:0]  io_out_memAddr,
  output         io_out_rdEn,
  output [4:0]   io_out_rdAddr,
  output [63:0]  io_out_rs1Data,
  output [63:0]  io_out_rs2Data,
  output [63:0]  io_out_imm,
  output [63:0]  io_out_aluRes,
  output [63:0]  io_out_memData,
  output [3:0]   io_out_csrOp,
  output         io_out_takenPre,
  output [31:0]  io_out_takenPrePC,
  output [63:0]  io_memRdData,
  output         io_memDone,
  output         io_memX1En,
  output [63:0]  io_memAluRes,
  output         io_cmp_ren,
  output         io_cmp_wen,
  output [63:0]  io_cmp_addr,
  output [63:0]  io_cmp_wdata,
  input  [63:0]  io_cmp_rdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire [63:0] _GEN_4 = io_in_aluRes % 64'h10; // @[DataMem.scala 37:27]
  wire [4:0] alignBits = _GEN_4[4:0]; // @[DataMem.scala 37:27]
  wire  _cmpWEn_T_3 = io_in_aluRes == 64'h2004000 | io_in_aluRes == 64'h200bff8; // @[DataMem.scala 40:59]
  wire  cmpWEn = io_in_memWr & (io_in_aluRes == 64'h2004000 | io_in_aluRes == 64'h200bff8); // @[DataMem.scala 40:32]
  wire  _cmpREn_T = io_in_memtoReg == 2'h1; // @[DataMem.scala 41:26]
  wire  cmpREn = io_in_memtoReg == 2'h1 & _cmpWEn_T_3; // @[DataMem.scala 41:35]
  wire  _dmemEn_T_6 = _cmpREn_T | io_in_memWr; // @[DataMem.scala 43:43]
  wire  dmemEn = ~(io_in_aluRes < 64'h80000000 | io_in_aluRes > 64'h88000000) & _dmemEn_T_6; // @[DataMem.scala 42:74]
  reg  dmemDone; // @[DataMem.scala 46:25]
  reg [31:0] inst; // @[DataMem.scala 47:17]
  wire  _T_2 = inst != io_in_inst; // @[DataMem.scala 52:54]
  wire  _GEN_0 = io_dmem_data_valid & io_IFDone & inst != io_in_inst ? 1'h0 : dmemDone; // @[DataMem.scala 52:70 53:14 46:25]
  wire  _GEN_1 = io_dmem_data_ready & io_IFDone | _GEN_0; // @[DataMem.scala 50:41 51:14]
  wire [63:0] _io_dmem_data_addr_T = io_dmem_data_valid ? io_in_aluRes : 64'h0; // @[DataMem.scala 61:27]
  wire [8:0] _io_dmem_data_write_T = alignBits * 4'h8; // @[DataMem.scala 62:48]
  wire [574:0] _GEN_5 = {{511'd0}, io_in_rs2Data}; // @[DataMem.scala 62:35]
  wire [574:0] _io_dmem_data_write_T_1 = _GEN_5 << _io_dmem_data_write_T; // @[DataMem.scala 62:35]
  wire [1:0] _io_dmem_data_strb_T_1 = 5'h1 == alignBits ? 2'h2 : 2'h1; // @[Mux.scala 81:58]
  wire [2:0] _io_dmem_data_strb_T_3 = 5'h2 == alignBits ? 3'h4 : {{1'd0}, _io_dmem_data_strb_T_1}; // @[Mux.scala 81:58]
  wire [3:0] _io_dmem_data_strb_T_5 = 5'h3 == alignBits ? 4'h8 : {{1'd0}, _io_dmem_data_strb_T_3}; // @[Mux.scala 81:58]
  wire [4:0] _io_dmem_data_strb_T_7 = 5'h4 == alignBits ? 5'h10 : {{1'd0}, _io_dmem_data_strb_T_5}; // @[Mux.scala 81:58]
  wire [5:0] _io_dmem_data_strb_T_9 = 5'h5 == alignBits ? 6'h20 : {{1'd0}, _io_dmem_data_strb_T_7}; // @[Mux.scala 81:58]
  wire [6:0] _io_dmem_data_strb_T_11 = 5'h6 == alignBits ? 7'h40 : {{1'd0}, _io_dmem_data_strb_T_9}; // @[Mux.scala 81:58]
  wire [7:0] _io_dmem_data_strb_T_13 = 5'h7 == alignBits ? 8'h80 : {{1'd0}, _io_dmem_data_strb_T_11}; // @[Mux.scala 81:58]
  wire [7:0] _io_dmem_data_strb_T_15 = 5'h9 == alignBits ? 8'h2 : _io_dmem_data_strb_T_13; // @[Mux.scala 81:58]
  wire [7:0] _io_dmem_data_strb_T_17 = 5'ha == alignBits ? 8'h4 : _io_dmem_data_strb_T_15; // @[Mux.scala 81:58]
  wire [7:0] _io_dmem_data_strb_T_19 = 5'hb == alignBits ? 8'h8 : _io_dmem_data_strb_T_17; // @[Mux.scala 81:58]
  wire [7:0] _io_dmem_data_strb_T_21 = 5'hc == alignBits ? 8'h10 : _io_dmem_data_strb_T_19; // @[Mux.scala 81:58]
  wire [7:0] _io_dmem_data_strb_T_23 = 5'hd == alignBits ? 8'h20 : _io_dmem_data_strb_T_21; // @[Mux.scala 81:58]
  wire [7:0] _io_dmem_data_strb_T_25 = 5'he == alignBits ? 8'h40 : _io_dmem_data_strb_T_23; // @[Mux.scala 81:58]
  wire [7:0] _io_dmem_data_strb_T_27 = 5'hf == alignBits ? 8'h80 : _io_dmem_data_strb_T_25; // @[Mux.scala 81:58]
  wire [3:0] _io_dmem_data_strb_T_29 = 5'h2 == alignBits ? 4'hc : 4'h3; // @[Mux.scala 81:58]
  wire [5:0] _io_dmem_data_strb_T_31 = 5'h4 == alignBits ? 6'h30 : {{2'd0}, _io_dmem_data_strb_T_29}; // @[Mux.scala 81:58]
  wire [7:0] _io_dmem_data_strb_T_33 = 5'h6 == alignBits ? 8'hc0 : {{2'd0}, _io_dmem_data_strb_T_31}; // @[Mux.scala 81:58]
  wire [7:0] _io_dmem_data_strb_T_35 = 5'ha == alignBits ? 8'hc : _io_dmem_data_strb_T_33; // @[Mux.scala 81:58]
  wire [7:0] _io_dmem_data_strb_T_37 = 5'hc == alignBits ? 8'h30 : _io_dmem_data_strb_T_35; // @[Mux.scala 81:58]
  wire [7:0] _io_dmem_data_strb_T_39 = 5'he == alignBits ? 8'hc0 : _io_dmem_data_strb_T_37; // @[Mux.scala 81:58]
  wire [7:0] _io_dmem_data_strb_T_43 = alignBits == 5'h0 | alignBits == 5'h8 ? 8'hf : 8'hf0; // @[DataMem.scala 92:22]
  wire [7:0] _io_dmem_data_strb_T_45 = 3'h0 == io_in_memOp ? _io_dmem_data_strb_T_27 : 8'h0; // @[Mux.scala 81:58]
  wire [7:0] _io_dmem_data_strb_T_47 = 3'h1 == io_in_memOp ? _io_dmem_data_strb_T_39 : _io_dmem_data_strb_T_45; // @[Mux.scala 81:58]
  wire [7:0] _io_dmem_data_strb_T_49 = 3'h2 == io_in_memOp ? _io_dmem_data_strb_T_43 : _io_dmem_data_strb_T_47; // @[Mux.scala 81:58]
  wire [7:0] _io_dmem_data_strb_T_51 = 3'h3 == io_in_memOp ? 8'hff : _io_dmem_data_strb_T_49; // @[Mux.scala 81:58]
  wire  dmemFire = io_dmem_data_valid & io_dmem_data_ready; // @[DataMem.scala 97:37]
  reg [63:0] rdata; // @[DataMem.scala 98:22]
  wire  _io_memDone_T_3 = _T_2 & dmemEn ? 1'h0 : dmemDone; // @[DataMem.scala 106:22]
  wire  rData_signBit = rdata[7]; // @[BitUtils.scala 18:20]
  wire [55:0] _rData_T_2 = rData_signBit ? 56'hffffffffffffff : 56'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _rData_T_3 = {_rData_T_2,rdata[7:0]}; // @[Cat.scala 31:58]
  wire  rData_signBit_1 = rdata[15]; // @[BitUtils.scala 18:20]
  wire [47:0] _rData_T_6 = rData_signBit_1 ? 48'hffffffffffff : 48'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _rData_T_7 = {_rData_T_6,rdata[15:0]}; // @[Cat.scala 31:58]
  wire  rData_signBit_2 = rdata[31]; // @[BitUtils.scala 18:20]
  wire [31:0] _rData_T_10 = rData_signBit_2 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _rData_T_11 = {_rData_T_10,rdata[31:0]}; // @[Cat.scala 31:58]
  wire [63:0] _rData_T_13 = {56'h0,rdata[7:0]}; // @[Cat.scala 31:58]
  wire [63:0] _rData_T_15 = {48'h0,rdata[15:0]}; // @[Cat.scala 31:58]
  wire [63:0] _rData_T_17 = {32'h0,rdata[31:0]}; // @[Cat.scala 31:58]
  wire [63:0] _rData_T_19 = 3'h0 == io_in_memOp ? _rData_T_3 : 64'h0; // @[Mux.scala 81:58]
  wire [63:0] _rData_T_21 = 3'h1 == io_in_memOp ? _rData_T_7 : _rData_T_19; // @[Mux.scala 81:58]
  wire [63:0] _rData_T_23 = 3'h2 == io_in_memOp ? _rData_T_11 : _rData_T_21; // @[Mux.scala 81:58]
  wire [63:0] _rData_T_25 = 3'h3 == io_in_memOp ? rdata : _rData_T_23; // @[Mux.scala 81:58]
  wire [63:0] _rData_T_27 = 3'h4 == io_in_memOp ? _rData_T_13 : _rData_T_25; // @[Mux.scala 81:58]
  wire [63:0] _rData_T_29 = 3'h5 == io_in_memOp ? _rData_T_15 : _rData_T_27; // @[Mux.scala 81:58]
  wire [63:0] rData = 3'h6 == io_in_memOp ? _rData_T_17 : _rData_T_29; // @[Mux.scala 81:58]
  wire  _data_size_T_7 = 3'h5 == io_in_memOp | 3'h1 == io_in_memOp; // @[Mux.scala 81:58]
  wire [1:0] _data_size_T_9 = 3'h3 == io_in_memOp ? 2'h3 : {{1'd0}, _data_size_T_7}; // @[Mux.scala 81:58]
  wire [1:0] _data_size_T_11 = 3'h2 == io_in_memOp ? 2'h2 : _data_size_T_9; // @[Mux.scala 81:58]
  wire [63:0] memData = io_in_memWr ? 64'h0 : rData; // @[DataMem.scala 159:18]
  wire  resW_signBit = io_in_aluRes[31]; // @[BitUtils.scala 18:20]
  wire [31:0] _resW_T_2 = resW_signBit ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] resW = {_resW_T_2,io_in_aluRes[31:0]}; // @[Cat.scala 31:58]
  wire [63:0] _memBPData_T_1 = 2'h0 == io_in_memtoReg ? io_in_aluRes : 64'h0; // @[Mux.scala 81:58]
  wire [63:0] _memBPData_T_3 = 2'h1 == io_in_memtoReg ? memData : _memBPData_T_1; // @[Mux.scala 81:58]
  wire [127:0] _io_cmp_wdata_T = cmpWEn ? io_dmem_data_write : 128'h0; // @[DataMem.scala 172:22]
  assign io_dmem_data_valid = ~io_memDone; // @[DataMem.scala 60:25]
  assign io_dmem_data_req = io_in_memWr & ~cmpWEn; // @[DataMem.scala 63:41]
  assign io_dmem_data_addr = _io_dmem_data_addr_T[31:0]; // @[DataMem.scala 61:21]
  assign io_dmem_data_size = 3'h6 == io_in_memOp ? 2'h2 : _data_size_T_11; // @[Mux.scala 81:58]
  assign io_dmem_data_strb = io_in_typeL ? 8'h0 : _io_dmem_data_strb_T_51; // @[DataMem.scala 65:27]
  assign io_dmem_data_write = _io_dmem_data_write_T_1[127:0]; // @[DataMem.scala 62:22]
  assign io_out_valid = io_in_valid; // @[DataMem.scala 200:19]
  assign io_out_pc = io_in_pc; // @[DataMem.scala 201:19]
  assign io_out_inst = io_in_inst; // @[DataMem.scala 202:19]
  assign io_out_typeL = io_in_typeL; // @[DataMem.scala 203:19]
  assign io_out_aluA = io_in_aluA; // @[DataMem.scala 204:19]
  assign io_out_aluB = io_in_aluB; // @[DataMem.scala 205:19]
  assign io_out_aluOp = io_in_aluOp; // @[DataMem.scala 206:19]
  assign io_out_branch = io_in_branch; // @[DataMem.scala 207:19]
  assign io_out_memtoReg = io_in_memtoReg; // @[DataMem.scala 208:19]
  assign io_out_memWr = io_in_memWr; // @[DataMem.scala 209:19]
  assign io_out_memOp = io_in_memOp; // @[DataMem.scala 210:19]
  assign io_out_memAddr = io_in_aluRes[31:0]; // @[DataMem.scala 211:19]
  assign io_out_rdEn = io_in_rdEn; // @[DataMem.scala 212:19]
  assign io_out_rdAddr = io_in_rdAddr; // @[DataMem.scala 213:19]
  assign io_out_rs1Data = io_in_rs1Data; // @[DataMem.scala 214:19]
  assign io_out_rs2Data = io_in_rs2Data; // @[DataMem.scala 215:19]
  assign io_out_imm = io_in_imm; // @[DataMem.scala 216:19]
  assign io_out_aluRes = io_in_aluRes; // @[DataMem.scala 219:19]
  assign io_out_memData = io_in_memWr ? 64'h0 : rData; // @[DataMem.scala 159:18]
  assign io_out_csrOp = io_in_csrOp; // @[DataMem.scala 221:19]
  assign io_out_takenPre = io_in_takenPre; // @[DataMem.scala 222:19]
  assign io_out_takenPrePC = io_in_takenPrePC; // @[DataMem.scala 223:21]
  assign io_memRdData = 2'h2 == io_in_memtoReg ? resW : _memBPData_T_3; // @[Mux.scala 81:58]
  assign io_memDone = cmpREn | cmpWEn | _io_memDone_T_3; // @[DataMem.scala 105:20]
  assign io_memX1En = io_in_rdEn & io_in_rdAddr == 5'h1; // @[DataMem.scala 228:28]
  assign io_memAluRes = io_in_aluRes; // @[DataMem.scala 229:16]
  assign io_cmp_ren = io_in_memtoReg == 2'h1 & _cmpWEn_T_3; // @[DataMem.scala 41:35]
  assign io_cmp_wen = io_in_memWr & (io_in_aluRes == 64'h2004000 | io_in_aluRes == 64'h200bff8); // @[DataMem.scala 40:32]
  assign io_cmp_addr = io_in_aluRes; // @[DataMem.scala 171:15]
  assign io_cmp_wdata = _io_cmp_wdata_T[63:0]; // @[DataMem.scala 172:16]
  always @(posedge clock) begin
    dmemDone <= reset | _GEN_1; // @[DataMem.scala 46:{25,25}]
    inst <= io_in_inst; // @[DataMem.scala 48:8]
    if (reset) begin // @[DataMem.scala 98:22]
      rdata <= 64'h0; // @[DataMem.scala 98:22]
    end else if (dmemFire) begin // @[DataMem.scala 99:18]
      rdata <= io_dmem_data_read; // @[DataMem.scala 100:11]
    end else if (cmpREn) begin // @[DataMem.scala 101:24]
      rdata <= io_cmp_rdata; // @[DataMem.scala 102:11]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  dmemDone = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  inst = _RAND_1[31:0];
  _RAND_2 = {2{`RANDOM}};
  rdata = _RAND_2[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CSR(
  input         clock,
  input         reset,
  input  [31:0] io_pc,
  input  [31:0] io_inst,
  input         io_csrEn,
  input  [63:0] io_rs1Data,
  input  [3:0]  io_csrOp,
  input  [11:0] io_rAddr,
  input         io_intr,
  output [63:0] io_rData,
  output [63:0] io_mepc,
  output [63:0] io_mtvec,
  output [63:0] io_mie,
  output [63:0] io_mstatus
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
`endif // RANDOMIZE_REG_INIT
  wire  dt_cs_clock; // @[CSR.scala 137:21]
  wire [7:0] dt_cs_coreid; // @[CSR.scala 137:21]
  wire [1:0] dt_cs_priviledgeMode; // @[CSR.scala 137:21]
  wire [63:0] dt_cs_mstatus; // @[CSR.scala 137:21]
  wire [63:0] dt_cs_sstatus; // @[CSR.scala 137:21]
  wire [63:0] dt_cs_mepc; // @[CSR.scala 137:21]
  wire [63:0] dt_cs_sepc; // @[CSR.scala 137:21]
  wire [63:0] dt_cs_mtval; // @[CSR.scala 137:21]
  wire [63:0] dt_cs_stval; // @[CSR.scala 137:21]
  wire [63:0] dt_cs_mtvec; // @[CSR.scala 137:21]
  wire [63:0] dt_cs_stvec; // @[CSR.scala 137:21]
  wire [63:0] dt_cs_mcause; // @[CSR.scala 137:21]
  wire [63:0] dt_cs_scause; // @[CSR.scala 137:21]
  wire [63:0] dt_cs_satp; // @[CSR.scala 137:21]
  wire [63:0] dt_cs_mip; // @[CSR.scala 137:21]
  wire [63:0] dt_cs_mie; // @[CSR.scala 137:21]
  wire [63:0] dt_cs_mscratch; // @[CSR.scala 137:21]
  wire [63:0] dt_cs_sscratch; // @[CSR.scala 137:21]
  wire [63:0] dt_cs_mideleg; // @[CSR.scala 137:21]
  wire [63:0] dt_cs_medeleg; // @[CSR.scala 137:21]
  reg [63:0] mstatus; // @[CSR.scala 29:24]
  reg [63:0] mtvec; // @[CSR.scala 30:24]
  reg [63:0] mepc; // @[CSR.scala 31:24]
  reg [63:0] mcause; // @[CSR.scala 32:24]
  reg [63:0] mie; // @[CSR.scala 35:26]
  reg [63:0] mscratch; // @[CSR.scala 37:26]
  reg [63:0] mcycle; // @[CSR.scala 38:26]
  wire [11:0] wAddr = io_inst[31:20]; // @[CSR.scala 49:24]
  wire [63:0] _rs1Data_T_3 = {59'h0,io_inst[19:15]}; // @[Cat.scala 31:58]
  wire [63:0] rs1Data = io_csrOp[2] ? _rs1Data_T_3 : io_rs1Data; // @[CSR.scala 52:20]
  wire  csrRW = ~io_csrOp[3] & io_csrOp != 4'h0; // @[CSR.scala 55:35]
  wire [63:0] _op1_T_1 = 12'h300 == wAddr ? mstatus : 64'h0; // @[Mux.scala 81:58]
  wire [63:0] _op1_T_3 = 12'h342 == wAddr ? mcause : _op1_T_1; // @[Mux.scala 81:58]
  wire [63:0] _op1_T_5 = 12'h304 == wAddr ? mie : _op1_T_3; // @[Mux.scala 81:58]
  wire [63:0] _op1_T_7 = 12'h305 == wAddr ? mtvec : _op1_T_5; // @[Mux.scala 81:58]
  wire [63:0] _op1_T_9 = 12'h340 == wAddr ? mscratch : _op1_T_7; // @[Mux.scala 81:58]
  wire [63:0] _op1_T_11 = 12'h341 == wAddr ? mepc : _op1_T_9; // @[Mux.scala 81:58]
  wire [63:0] _op1_T_13 = 12'h344 == wAddr ? 64'h0 : _op1_T_11; // @[Mux.scala 81:58]
  wire [63:0] _op1_T_15 = 12'hb00 == wAddr ? mcycle : _op1_T_13; // @[Mux.scala 81:58]
  wire [63:0] op1 = 12'hb02 == wAddr ? 64'h0 : _op1_T_15; // @[Mux.scala 81:58]
  wire [63:0] _wdata_T_1 = op1 | rs1Data; // @[CSR.scala 71:23]
  wire [63:0] _wdata_T_2 = ~rs1Data; // @[CSR.scala 72:25]
  wire [63:0] _wdata_T_3 = op1 & _wdata_T_2; // @[CSR.scala 72:23]
  wire [63:0] _wdata_T_5 = 2'h1 == io_csrOp[1:0] ? rs1Data : 64'h0; // @[Mux.scala 81:58]
  wire [63:0] _wdata_T_7 = 2'h2 == io_csrOp[1:0] ? _wdata_T_1 : _wdata_T_5; // @[Mux.scala 81:58]
  wire [63:0] _wdata_T_9 = 2'h3 == io_csrOp[1:0] ? _wdata_T_3 : _wdata_T_7; // @[Mux.scala 81:58]
  wire [63:0] wdata = csrRW ? _wdata_T_9 : 64'h0; // @[CSR.scala 68:18]
  wire [63:0] _mstatus_T_5 = {mstatus[63:13],2'h3,mstatus[10:8],mstatus[3],mstatus[6:4],1'h0,mstatus[2:0]}; // @[Cat.scala 31:58]
  wire [63:0] _mstatus_T_11 = {mstatus[63:13],2'h0,mstatus[10:8],1'h1,mstatus[6:4],mstatus[7],mstatus[2:0]}; // @[Cat.scala 31:58]
  wire [63:0] _GEN_0 = io_intr & io_csrEn ? {{32'd0}, io_pc} : mepc; // @[CSR.scala 85:33 87:10 31:24]
  wire [63:0] _GEN_1 = io_intr & io_csrEn ? 64'h8000000000000007 : mcause; // @[CSR.scala 85:33 88:12 32:24]
  wire [63:0] _GEN_2 = io_intr & io_csrEn ? _mstatus_T_5 : mstatus; // @[CSR.scala 85:33 89:13 29:24]
  wire [63:0] _GEN_3 = io_csrOp == 4'h9 & io_csrEn ? _mstatus_T_11 : _GEN_2; // @[CSR.scala 82:50 84:13]
  wire [63:0] _GEN_4 = io_csrOp == 4'h9 & io_csrEn ? mepc : _GEN_0; // @[CSR.scala 31:24 82:50]
  wire [63:0] _GEN_5 = io_csrOp == 4'h9 & io_csrEn ? mcause : _GEN_1; // @[CSR.scala 32:24 82:50]
  wire [63:0] _GEN_6 = io_csrOp == 4'h8 & io_csrEn ? 64'hb : _GEN_5; // @[CSR.scala 77:43 79:13]
  wire [63:0] _GEN_7 = io_csrOp == 4'h8 & io_csrEn ? {{32'd0}, io_pc} : _GEN_4; // @[CSR.scala 77:43 80:13]
  wire [63:0] _GEN_8 = io_csrOp == 4'h8 & io_csrEn ? _mstatus_T_5 : _GEN_3; // @[CSR.scala 77:43 81:13]
  reg [63:0] mtvec_REG; // @[CSR.scala 99:23]
  wire  _mstatus_T_24 = wdata[16] & wdata[15] | wdata[14] & wdata[13]; // @[CSR.scala 108:46]
  wire [63:0] _mstatus_T_26 = {_mstatus_T_24,wdata[62:0]}; // @[Cat.scala 31:58]
  reg [63:0] mie_REG; // @[CSR.scala 111:21]
  wire [63:0] _io_rData_T_1 = 12'h300 == io_rAddr ? mstatus : 64'h0; // @[Mux.scala 81:58]
  wire [63:0] _io_rData_T_3 = 12'h342 == io_rAddr ? mcause : _io_rData_T_1; // @[Mux.scala 81:58]
  wire [63:0] _io_rData_T_5 = 12'h304 == io_rAddr ? mie : _io_rData_T_3; // @[Mux.scala 81:58]
  wire [63:0] _io_rData_T_7 = 12'h305 == io_rAddr ? mtvec : _io_rData_T_5; // @[Mux.scala 81:58]
  wire [63:0] _io_rData_T_9 = 12'h340 == io_rAddr ? mscratch : _io_rData_T_7; // @[Mux.scala 81:58]
  wire [63:0] _io_rData_T_11 = 12'h341 == io_rAddr ? mepc : _io_rData_T_9; // @[Mux.scala 81:58]
  wire [63:0] _io_rData_T_13 = 12'h344 == io_rAddr ? 64'h0 : _io_rData_T_11; // @[Mux.scala 81:58]
  wire [63:0] _io_rData_T_15 = 12'hb00 == io_rAddr ? mcycle : _io_rData_T_13; // @[Mux.scala 81:58]
  DifftestCSRState dt_cs ( // @[CSR.scala 137:21]
    .clock(dt_cs_clock),
    .coreid(dt_cs_coreid),
    .priviledgeMode(dt_cs_priviledgeMode),
    .mstatus(dt_cs_mstatus),
    .sstatus(dt_cs_sstatus),
    .mepc(dt_cs_mepc),
    .sepc(dt_cs_sepc),
    .mtval(dt_cs_mtval),
    .stval(dt_cs_stval),
    .mtvec(dt_cs_mtvec),
    .stvec(dt_cs_stvec),
    .mcause(dt_cs_mcause),
    .scause(dt_cs_scause),
    .satp(dt_cs_satp),
    .mip(dt_cs_mip),
    .mie(dt_cs_mie),
    .mscratch(dt_cs_mscratch),
    .sscratch(dt_cs_sscratch),
    .mideleg(dt_cs_mideleg),
    .medeleg(dt_cs_medeleg)
  );
  assign io_rData = 12'hb02 == io_rAddr ? 64'h0 : _io_rData_T_15; // @[Mux.scala 81:58]
  assign io_mepc = mepc; // @[CSR.scala 131:11]
  assign io_mtvec = mtvec; // @[CSR.scala 132:12]
  assign io_mie = mie; // @[CSR.scala 133:10]
  assign io_mstatus = mstatus; // @[CSR.scala 134:14]
  assign dt_cs_clock = clock; // @[CSR.scala 138:27]
  assign dt_cs_coreid = 8'h0; // @[CSR.scala 139:27]
  assign dt_cs_priviledgeMode = 2'h3; // @[CSR.scala 140:27]
  assign dt_cs_mstatus = mstatus; // @[CSR.scala 141:27]
  assign dt_cs_sstatus = mstatus & 64'h80000003000de122; // @[CSR.scala 142:38]
  assign dt_cs_mepc = mepc; // @[CSR.scala 143:27]
  assign dt_cs_sepc = 64'h0; // @[CSR.scala 144:27]
  assign dt_cs_mtval = 64'h0; // @[CSR.scala 145:27]
  assign dt_cs_stval = 64'h0; // @[CSR.scala 146:27]
  assign dt_cs_mtvec = mtvec; // @[CSR.scala 147:27]
  assign dt_cs_stvec = 64'h0; // @[CSR.scala 148:27]
  assign dt_cs_mcause = mcause; // @[CSR.scala 149:27]
  assign dt_cs_scause = 64'h0; // @[CSR.scala 150:27]
  assign dt_cs_satp = 64'h0; // @[CSR.scala 151:27]
  assign dt_cs_mip = 64'h0; // @[CSR.scala 152:27]
  assign dt_cs_mie = mie; // @[CSR.scala 153:27]
  assign dt_cs_mscratch = mscratch; // @[CSR.scala 154:27]
  assign dt_cs_sscratch = 64'h0; // @[CSR.scala 155:27]
  assign dt_cs_mideleg = 64'h0; // @[CSR.scala 156:27]
  assign dt_cs_medeleg = 64'h0; // @[CSR.scala 157:27]
  always @(posedge clock) begin
    if (reset) begin // @[CSR.scala 29:24]
      mstatus <= 64'h1800; // @[CSR.scala 29:24]
    end else if (csrRW & io_csrEn & ~io_intr) begin // @[CSR.scala 94:36]
      if (wAddr == 12'h300) begin // @[CSR.scala 107:34]
        mstatus <= _mstatus_T_26; // @[CSR.scala 108:15]
      end else begin
        mstatus <= _GEN_8;
      end
    end else begin
      mstatus <= _GEN_8;
    end
    if (reset) begin // @[CSR.scala 30:24]
      mtvec <= 64'h0; // @[CSR.scala 30:24]
    end else if (csrRW & io_csrEn & ~io_intr) begin // @[CSR.scala 94:36]
      if (wAddr == 12'h305) begin // @[CSR.scala 98:32]
        mtvec <= mtvec_REG; // @[CSR.scala 99:13]
      end
    end
    if (reset) begin // @[CSR.scala 31:24]
      mepc <= 64'h0; // @[CSR.scala 31:24]
    end else if (csrRW & io_csrEn & ~io_intr) begin // @[CSR.scala 94:36]
      if (wAddr == 12'h341) begin // @[CSR.scala 101:31]
        if (csrRW) begin // @[CSR.scala 68:18]
          mepc <= _wdata_T_9;
        end else begin
          mepc <= 64'h0;
        end
      end else begin
        mepc <= _GEN_7;
      end
    end else begin
      mepc <= _GEN_7;
    end
    if (reset) begin // @[CSR.scala 32:24]
      mcause <= 64'h0; // @[CSR.scala 32:24]
    end else if (csrRW & io_csrEn & ~io_intr) begin // @[CSR.scala 94:36]
      if (wAddr == 12'h342) begin // @[CSR.scala 104:33]
        if (csrRW) begin // @[CSR.scala 68:18]
          mcause <= _wdata_T_9;
        end else begin
          mcause <= 64'h0;
        end
      end else begin
        mcause <= _GEN_6;
      end
    end else begin
      mcause <= _GEN_6;
    end
    if (reset) begin // @[CSR.scala 35:26]
      mie <= 64'h0; // @[CSR.scala 35:26]
    end else if (csrRW & io_csrEn & ~io_intr) begin // @[CSR.scala 94:36]
      if (wAddr == 12'h304) begin // @[CSR.scala 110:30]
        mie <= mie_REG; // @[CSR.scala 111:11]
      end
    end
    if (reset) begin // @[CSR.scala 37:26]
      mscratch <= 64'h0; // @[CSR.scala 37:26]
    end else if (csrRW & io_csrEn & ~io_intr) begin // @[CSR.scala 94:36]
      if (wAddr == 12'h340) begin // @[CSR.scala 113:35]
        if (csrRW) begin // @[CSR.scala 68:18]
          mscratch <= _wdata_T_9;
        end else begin
          mscratch <= 64'h0;
        end
      end
    end
    if (reset) begin // @[CSR.scala 38:26]
      mcycle <= 64'h0; // @[CSR.scala 38:26]
    end else if (csrRW & io_csrEn & ~io_intr) begin // @[CSR.scala 94:36]
      if (wAddr == 12'hb00) begin // @[CSR.scala 95:33]
        if (csrRW) begin // @[CSR.scala 68:18]
          mcycle <= _wdata_T_9;
        end else begin
          mcycle <= 64'h0;
        end
      end
    end
    if (csrRW) begin // @[CSR.scala 68:18]
      if (2'h3 == io_csrOp[1:0]) begin // @[Mux.scala 81:58]
        mtvec_REG <= _wdata_T_3;
      end else if (2'h2 == io_csrOp[1:0]) begin // @[Mux.scala 81:58]
        mtvec_REG <= _wdata_T_1;
      end else if (2'h1 == io_csrOp[1:0]) begin // @[Mux.scala 81:58]
        mtvec_REG <= rs1Data;
      end else begin
        mtvec_REG <= 64'h0;
      end
    end else begin
      mtvec_REG <= 64'h0;
    end
    if (csrRW) begin // @[CSR.scala 68:18]
      if (2'h3 == io_csrOp[1:0]) begin // @[Mux.scala 81:58]
        mie_REG <= _wdata_T_3;
      end else if (2'h2 == io_csrOp[1:0]) begin // @[Mux.scala 81:58]
        mie_REG <= _wdata_T_1;
      end else if (2'h1 == io_csrOp[1:0]) begin // @[Mux.scala 81:58]
        mie_REG <= rs1Data;
      end else begin
        mie_REG <= 64'h0;
      end
    end else begin
      mie_REG <= 64'h0;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  mstatus = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  mtvec = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  mepc = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  mcause = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  mie = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  mscratch = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  mcycle = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  mtvec_REG = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  mie_REG = _RAND_8[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CLINT(
  input         clock,
  input         reset,
  input  [63:0] io_mstatus,
  input  [63:0] io_mie,
  input         io_csrEn,
  input         io_cmp_ren,
  input         io_cmp_wen,
  input  [63:0] io_cmp_addr,
  input  [63:0] io_cmp_wdata,
  output [63:0] io_cmp_rdata,
  output        io_time_int
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] mtime; // @[CLINT.scala 22:22]
  reg [63:0] mtimecmp; // @[CLINT.scala 23:25]
  wire [63:0] _mtime_T_1 = mtime + 64'h1; // @[CLINT.scala 25:18]
  wire  _io_time_int_T_5 = mtime >= mtimecmp; // @[CLINT.scala 30:26]
  wire  _io_time_int_T_6 = io_mstatus[3] & io_mie[7] & _io_time_int_T_5; // @[CLINT.scala 29:64]
  wire [63:0] _io_cmp_rdata_T_1 = io_cmp_addr == 64'h200bff8 ? mtime : mtimecmp; // @[CLINT.scala 32:24]
  assign io_cmp_rdata = io_cmp_ren ? _io_cmp_rdata_T_1 : 64'h0; // @[CLINT.scala 31:22]
  assign io_time_int = _io_time_int_T_6 & io_csrEn; // @[CLINT.scala 30:40]
  always @(posedge clock) begin
    if (reset) begin // @[CLINT.scala 22:22]
      mtime <= 64'h0; // @[CLINT.scala 22:22]
    end else begin
      mtime <= _mtime_T_1; // @[CLINT.scala 25:9]
    end
    if (reset) begin // @[CLINT.scala 23:25]
      mtimecmp <= 64'h0; // @[CLINT.scala 23:25]
    end else if (io_cmp_wen) begin // @[CLINT.scala 26:21]
      mtimecmp <= io_cmp_wdata; // @[CLINT.scala 27:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  mtime = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  mtimecmp = _RAND_1[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module WriteBack(
  input         clock,
  input         reset,
  input         io_in_valid,
  input  [31:0] io_in_pc,
  input  [31:0] io_in_inst,
  input  [1:0]  io_in_memtoReg,
  input         io_in_memWr,
  input  [31:0] io_in_memAddr,
  input         io_in_rdEn,
  input  [4:0]  io_in_rdAddr,
  input  [63:0] io_in_rs1Data,
  input  [63:0] io_in_aluRes,
  input  [63:0] io_in_memData,
  input  [3:0]  io_in_csrOp,
  input         io_IFDone,
  input         io_memDone,
  input  [31:0] io_pc_intr,
  output [31:0] io_pc,
  output [31:0] io_inst,
  output        io_wbRdEn,
  output [4:0]  io_wbRdAddr,
  output [63:0] io_wbRdData,
  output        io_ready_cmt,
  output [3:0]  io_csrOp_WB,
  output [63:0] io_mepc,
  output [63:0] io_mtvec,
  input         io_cmp_ren,
  input         io_cmp_wen,
  input  [63:0] io_cmp_addr,
  input  [63:0] io_cmp_wdata,
  output [63:0] io_cmp_rdata,
  output        io_exc,
  output [1:0]  io_memtoReg,
  output        io_memWr,
  output [31:0] io_mem_addr,
  output        io_time_int
);
  wire  csr_clock; // @[WriteBack.scala 41:21]
  wire  csr_reset; // @[WriteBack.scala 41:21]
  wire [31:0] csr_io_pc; // @[WriteBack.scala 41:21]
  wire [31:0] csr_io_inst; // @[WriteBack.scala 41:21]
  wire  csr_io_csrEn; // @[WriteBack.scala 41:21]
  wire [63:0] csr_io_rs1Data; // @[WriteBack.scala 41:21]
  wire [3:0] csr_io_csrOp; // @[WriteBack.scala 41:21]
  wire [11:0] csr_io_rAddr; // @[WriteBack.scala 41:21]
  wire  csr_io_intr; // @[WriteBack.scala 41:21]
  wire [63:0] csr_io_rData; // @[WriteBack.scala 41:21]
  wire [63:0] csr_io_mepc; // @[WriteBack.scala 41:21]
  wire [63:0] csr_io_mtvec; // @[WriteBack.scala 41:21]
  wire [63:0] csr_io_mie; // @[WriteBack.scala 41:21]
  wire [63:0] csr_io_mstatus; // @[WriteBack.scala 41:21]
  wire  clint_clock; // @[WriteBack.scala 42:23]
  wire  clint_reset; // @[WriteBack.scala 42:23]
  wire [63:0] clint_io_mstatus; // @[WriteBack.scala 42:23]
  wire [63:0] clint_io_mie; // @[WriteBack.scala 42:23]
  wire  clint_io_csrEn; // @[WriteBack.scala 42:23]
  wire  clint_io_cmp_ren; // @[WriteBack.scala 42:23]
  wire  clint_io_cmp_wen; // @[WriteBack.scala 42:23]
  wire [63:0] clint_io_cmp_addr; // @[WriteBack.scala 42:23]
  wire [63:0] clint_io_cmp_wdata; // @[WriteBack.scala 42:23]
  wire [63:0] clint_io_cmp_rdata; // @[WriteBack.scala 42:23]
  wire  clint_io_time_int; // @[WriteBack.scala 42:23]
  wire  csrEn = io_IFDone & io_memDone; // @[WriteBack.scala 44:27]
  wire  resW_signBit = io_in_aluRes[31]; // @[BitUtils.scala 18:20]
  wire [31:0] _resW_T_2 = resW_signBit ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] resW = {_resW_T_2,io_in_aluRes[31:0]}; // @[Cat.scala 31:58]
  wire [63:0] _rdData_T_1 = 2'h0 == io_in_memtoReg ? io_in_aluRes : 64'h0; // @[Mux.scala 81:58]
  wire [63:0] _rdData_T_3 = 2'h1 == io_in_memtoReg ? io_in_memData : _rdData_T_1; // @[Mux.scala 81:58]
  wire [63:0] rdData = 2'h2 == io_in_memtoReg ? resW : _rdData_T_3; // @[Mux.scala 81:58]
  wire [4:0] _io_wbRdAddr_T = clint_io_time_int ? 5'h0 : io_in_rdAddr; // @[WriteBack.scala 75:32]
  wire [63:0] _io_wbRdData_T_1 = io_in_csrOp == 4'h0 ? rdData : csr_io_rData; // @[WriteBack.scala 76:32]
  wire  _io_ready_cmt_T_1 = ~clint_io_time_int; // @[WriteBack.scala 79:21]
  wire  _io_ready_cmt_T_2 = io_in_inst != 32'h0 & _io_ready_cmt_T_1; // @[WriteBack.scala 78:38]
  wire  _io_ready_cmt_T_3 = csrEn ? io_IFDone : io_in_valid; // @[WriteBack.scala 80:27]
  CSR csr ( // @[WriteBack.scala 41:21]
    .clock(csr_clock),
    .reset(csr_reset),
    .io_pc(csr_io_pc),
    .io_inst(csr_io_inst),
    .io_csrEn(csr_io_csrEn),
    .io_rs1Data(csr_io_rs1Data),
    .io_csrOp(csr_io_csrOp),
    .io_rAddr(csr_io_rAddr),
    .io_intr(csr_io_intr),
    .io_rData(csr_io_rData),
    .io_mepc(csr_io_mepc),
    .io_mtvec(csr_io_mtvec),
    .io_mie(csr_io_mie),
    .io_mstatus(csr_io_mstatus)
  );
  CLINT clint ( // @[WriteBack.scala 42:23]
    .clock(clint_clock),
    .reset(clint_reset),
    .io_mstatus(clint_io_mstatus),
    .io_mie(clint_io_mie),
    .io_csrEn(clint_io_csrEn),
    .io_cmp_ren(clint_io_cmp_ren),
    .io_cmp_wen(clint_io_cmp_wen),
    .io_cmp_addr(clint_io_cmp_addr),
    .io_cmp_wdata(clint_io_cmp_wdata),
    .io_cmp_rdata(clint_io_cmp_rdata),
    .io_time_int(clint_io_time_int)
  );
  assign io_pc = io_in_pc; // @[WriteBack.scala 71:9]
  assign io_inst = io_in_inst; // @[WriteBack.scala 72:11]
  assign io_wbRdEn = csrEn & io_in_rdEn; // @[WriteBack.scala 74:19]
  assign io_wbRdAddr = csrEn ? _io_wbRdAddr_T : 5'h0; // @[WriteBack.scala 75:21]
  assign io_wbRdData = csrEn ? _io_wbRdData_T_1 : 64'h0; // @[WriteBack.scala 76:21]
  assign io_ready_cmt = _io_ready_cmt_T_2 & _io_ready_cmt_T_3; // @[WriteBack.scala 79:40]
  assign io_csrOp_WB = io_in_csrOp; // @[WriteBack.scala 84:15]
  assign io_mepc = csr_io_mepc; // @[WriteBack.scala 82:14]
  assign io_mtvec = csr_io_mtvec; // @[WriteBack.scala 83:14]
  assign io_cmp_rdata = clint_io_cmp_rdata; // @[WriteBack.scala 85:16]
  assign io_exc = io_in_csrOp[3] | clint_io_time_int; // @[WriteBack.scala 90:37]
  assign io_memtoReg = io_in_memtoReg; // @[WriteBack.scala 87:15]
  assign io_memWr = io_in_memWr; // @[WriteBack.scala 88:12]
  assign io_mem_addr = io_in_memAddr; // @[WriteBack.scala 89:15]
  assign io_time_int = clint_io_time_int; // @[WriteBack.scala 92:15]
  assign csr_clock = clock;
  assign csr_reset = reset;
  assign csr_io_pc = clint_io_time_int ? io_pc_intr : io_in_pc; // @[WriteBack.scala 46:21]
  assign csr_io_inst = io_in_inst; // @[WriteBack.scala 47:17]
  assign csr_io_csrEn = io_IFDone & io_memDone; // @[WriteBack.scala 44:27]
  assign csr_io_rs1Data = io_in_rs1Data; // @[WriteBack.scala 49:20]
  assign csr_io_csrOp = io_in_csrOp; // @[WriteBack.scala 50:18]
  assign csr_io_rAddr = io_in_inst[31:20]; // @[WriteBack.scala 51:31]
  assign csr_io_intr = clint_io_time_int; // @[WriteBack.scala 52:17]
  assign clint_clock = clock;
  assign clint_reset = reset;
  assign clint_io_mstatus = csr_io_mstatus; // @[WriteBack.scala 54:22]
  assign clint_io_mie = csr_io_mie; // @[WriteBack.scala 55:18]
  assign clint_io_csrEn = io_IFDone & io_memDone; // @[WriteBack.scala 44:27]
  assign clint_io_cmp_ren = io_cmp_ren; // @[WriteBack.scala 58:22]
  assign clint_io_cmp_wen = io_cmp_wen; // @[WriteBack.scala 59:22]
  assign clint_io_cmp_addr = io_cmp_addr; // @[WriteBack.scala 60:23]
  assign clint_io_cmp_wdata = io_cmp_wdata; // @[WriteBack.scala 61:24]
endmodule
module preDebug(
  input        clock,
  input        reset,
  input  [2:0] io_exeBranch,
  input        io_takenMiss,
  input  [4:0] io_rs1Addr,
  input        io_coreEnd,
  input        io_IFDone,
  input        io_memDone
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] bjp_0; // @[preDebug.scala 17:20]
  reg [31:0] bjp_1; // @[preDebug.scala 17:20]
  reg [31:0] bjp_2; // @[preDebug.scala 17:20]
  reg [31:0] bjp_3; // @[preDebug.scala 17:20]
  reg [31:0] bjp_4; // @[preDebug.scala 17:20]
  reg [31:0] bjp_5; // @[preDebug.scala 17:20]
  reg [31:0] bjp_6; // @[preDebug.scala 17:20]
  reg [31:0] bjpMiss_0; // @[preDebug.scala 18:24]
  reg [31:0] bjpMiss_1; // @[preDebug.scala 18:24]
  reg [31:0] bjpMiss_2; // @[preDebug.scala 18:24]
  reg [31:0] bjpMiss_3; // @[preDebug.scala 18:24]
  reg [31:0] bjpMiss_4; // @[preDebug.scala 18:24]
  reg [31:0] bjpMiss_5; // @[preDebug.scala 18:24]
  reg [31:0] bjpMiss_6; // @[preDebug.scala 18:24]
  wire [31:0] _bjp_0_T_1 = bjp_0 + 32'h1; // @[preDebug.scala 21:22]
  wire [31:0] _bjpMiss_0_T_1 = bjpMiss_0 + 32'h1; // @[preDebug.scala 23:32]
  wire [31:0] _bjp_6_T_1 = bjp_6 + 32'h1; // @[preDebug.scala 27:24]
  wire [31:0] _bjpMiss_6_T_1 = bjpMiss_6 + 32'h1; // @[preDebug.scala 29:34]
  wire [31:0] _GEN_1 = io_takenMiss ? _bjpMiss_6_T_1 : bjpMiss_6; // @[preDebug.scala 28:26 29:20 18:24]
  wire [31:0] _bjp_1_T_1 = bjp_1 + 32'h1; // @[preDebug.scala 32:24]
  wire [31:0] _bjpMiss_1_T_1 = bjpMiss_1 + 32'h1; // @[preDebug.scala 34:34]
  wire [31:0] _GEN_2 = io_takenMiss ? _bjpMiss_1_T_1 : bjpMiss_1; // @[preDebug.scala 33:26 34:20 18:24]
  wire [31:0] _GEN_3 = io_rs1Addr == 5'h1 ? _bjp_6_T_1 : bjp_6; // @[preDebug.scala 26:29 27:14 17:20]
  wire [31:0] _GEN_4 = io_rs1Addr == 5'h1 ? _GEN_1 : bjpMiss_6; // @[preDebug.scala 18:24 26:29]
  wire [31:0] _GEN_5 = io_rs1Addr == 5'h1 ? bjp_1 : _bjp_1_T_1; // @[preDebug.scala 17:20 26:29 32:14]
  wire [31:0] _GEN_6 = io_rs1Addr == 5'h1 ? bjpMiss_1 : _GEN_2; // @[preDebug.scala 18:24 26:29]
  wire [31:0] _bjp_2_T_1 = bjp_2 + 32'h1; // @[preDebug.scala 38:22]
  wire [31:0] _bjpMiss_2_T_1 = bjpMiss_2 + 32'h1; // @[preDebug.scala 40:32]
  wire [31:0] _GEN_7 = io_takenMiss ? _bjpMiss_2_T_1 : bjpMiss_2; // @[preDebug.scala 39:24 40:18 18:24]
  wire [31:0] _bjp_3_T_1 = bjp_3 + 32'h1; // @[preDebug.scala 43:22]
  wire [31:0] _bjpMiss_3_T_1 = bjpMiss_3 + 32'h1; // @[preDebug.scala 45:32]
  wire [31:0] _GEN_8 = io_takenMiss ? _bjpMiss_3_T_1 : bjpMiss_3; // @[preDebug.scala 44:24 45:18 18:24]
  wire [31:0] _bjp_4_T_1 = bjp_4 + 32'h1; // @[preDebug.scala 48:22]
  wire [31:0] _bjpMiss_4_T_1 = bjpMiss_4 + 32'h1; // @[preDebug.scala 50:32]
  wire [31:0] _GEN_9 = io_takenMiss ? _bjpMiss_4_T_1 : bjpMiss_4; // @[preDebug.scala 49:24 50:18 18:24]
  wire [31:0] _bjp_5_T_1 = bjp_5 + 32'h1; // @[preDebug.scala 53:22]
  wire [31:0] _bjpMiss_5_T_1 = bjpMiss_5 + 32'h1; // @[preDebug.scala 55:32]
  wire [31:0] _GEN_10 = io_takenMiss ? _bjpMiss_5_T_1 : bjpMiss_5; // @[preDebug.scala 54:24 55:18 18:24]
  wire [31:0] _GEN_11 = io_exeBranch == 3'h7 ? _bjp_5_T_1 : bjp_5; // @[preDebug.scala 52:43 53:12 17:20]
  wire [31:0] _GEN_12 = io_exeBranch == 3'h7 ? _GEN_10 : bjpMiss_5; // @[preDebug.scala 18:24 52:43]
  wire [31:0] _GEN_13 = io_exeBranch == 3'h6 ? _bjp_4_T_1 : bjp_4; // @[preDebug.scala 47:43 48:12 17:20]
  wire [31:0] _GEN_14 = io_exeBranch == 3'h6 ? _GEN_9 : bjpMiss_4; // @[preDebug.scala 18:24 47:43]
  wire [31:0] _GEN_15 = io_exeBranch == 3'h6 ? bjp_5 : _GEN_11; // @[preDebug.scala 17:20 47:43]
  wire [31:0] _GEN_16 = io_exeBranch == 3'h6 ? bjpMiss_5 : _GEN_12; // @[preDebug.scala 18:24 47:43]
  wire [31:0] _GEN_17 = io_exeBranch == 3'h5 ? _bjp_3_T_1 : bjp_3; // @[preDebug.scala 42:43 43:12 17:20]
  wire [31:0] _GEN_18 = io_exeBranch == 3'h5 ? _GEN_8 : bjpMiss_3; // @[preDebug.scala 18:24 42:43]
  wire [31:0] _GEN_19 = io_exeBranch == 3'h5 ? bjp_4 : _GEN_13; // @[preDebug.scala 17:20 42:43]
  wire [31:0] _GEN_20 = io_exeBranch == 3'h5 ? bjpMiss_4 : _GEN_14; // @[preDebug.scala 18:24 42:43]
  wire [31:0] _GEN_21 = io_exeBranch == 3'h5 ? bjp_5 : _GEN_15; // @[preDebug.scala 17:20 42:43]
  wire [31:0] _GEN_22 = io_exeBranch == 3'h5 ? bjpMiss_5 : _GEN_16; // @[preDebug.scala 18:24 42:43]
  wire [31:0] _GEN_23 = io_exeBranch == 3'h4 ? _bjp_2_T_1 : bjp_2; // @[preDebug.scala 37:43 38:12 17:20]
  wire [31:0] _GEN_24 = io_exeBranch == 3'h4 ? _GEN_7 : bjpMiss_2; // @[preDebug.scala 18:24 37:43]
  wire [31:0] _GEN_25 = io_exeBranch == 3'h4 ? bjp_3 : _GEN_17; // @[preDebug.scala 17:20 37:43]
  wire [31:0] _GEN_26 = io_exeBranch == 3'h4 ? bjpMiss_3 : _GEN_18; // @[preDebug.scala 18:24 37:43]
  wire [31:0] _GEN_27 = io_exeBranch == 3'h4 ? bjp_4 : _GEN_19; // @[preDebug.scala 17:20 37:43]
  wire [31:0] _GEN_28 = io_exeBranch == 3'h4 ? bjpMiss_4 : _GEN_20; // @[preDebug.scala 18:24 37:43]
  wire [31:0] _GEN_29 = io_exeBranch == 3'h4 ? bjp_5 : _GEN_21; // @[preDebug.scala 17:20 37:43]
  wire [31:0] _GEN_30 = io_exeBranch == 3'h4 ? bjpMiss_5 : _GEN_22; // @[preDebug.scala 18:24 37:43]
  wire  _T_9 = io_coreEnd & io_IFDone & io_memDone; // @[preDebug.scala 67:32]
  wire  _T_11 = ~reset; // @[preDebug.scala 68:11]
  always @(posedge clock) begin
    if (reset) begin // @[preDebug.scala 17:20]
      bjp_0 <= 32'h0; // @[preDebug.scala 17:20]
    end else if (io_IFDone & io_memDone) begin // @[preDebug.scala 19:31]
      if (io_exeBranch == 3'h1) begin // @[preDebug.scala 20:36]
        bjp_0 <= _bjp_0_T_1; // @[preDebug.scala 21:12]
      end
    end
    if (reset) begin // @[preDebug.scala 17:20]
      bjp_1 <= 32'h0; // @[preDebug.scala 17:20]
    end else if (io_IFDone & io_memDone) begin // @[preDebug.scala 19:31]
      if (!(io_exeBranch == 3'h1)) begin // @[preDebug.scala 20:36]
        if (io_exeBranch == 3'h2) begin // @[preDebug.scala 25:43]
          bjp_1 <= _GEN_5;
        end
      end
    end
    if (reset) begin // @[preDebug.scala 17:20]
      bjp_2 <= 32'h0; // @[preDebug.scala 17:20]
    end else if (io_IFDone & io_memDone) begin // @[preDebug.scala 19:31]
      if (!(io_exeBranch == 3'h1)) begin // @[preDebug.scala 20:36]
        if (!(io_exeBranch == 3'h2)) begin // @[preDebug.scala 25:43]
          bjp_2 <= _GEN_23;
        end
      end
    end
    if (reset) begin // @[preDebug.scala 17:20]
      bjp_3 <= 32'h0; // @[preDebug.scala 17:20]
    end else if (io_IFDone & io_memDone) begin // @[preDebug.scala 19:31]
      if (!(io_exeBranch == 3'h1)) begin // @[preDebug.scala 20:36]
        if (!(io_exeBranch == 3'h2)) begin // @[preDebug.scala 25:43]
          bjp_3 <= _GEN_25;
        end
      end
    end
    if (reset) begin // @[preDebug.scala 17:20]
      bjp_4 <= 32'h0; // @[preDebug.scala 17:20]
    end else if (io_IFDone & io_memDone) begin // @[preDebug.scala 19:31]
      if (!(io_exeBranch == 3'h1)) begin // @[preDebug.scala 20:36]
        if (!(io_exeBranch == 3'h2)) begin // @[preDebug.scala 25:43]
          bjp_4 <= _GEN_27;
        end
      end
    end
    if (reset) begin // @[preDebug.scala 17:20]
      bjp_5 <= 32'h0; // @[preDebug.scala 17:20]
    end else if (io_IFDone & io_memDone) begin // @[preDebug.scala 19:31]
      if (!(io_exeBranch == 3'h1)) begin // @[preDebug.scala 20:36]
        if (!(io_exeBranch == 3'h2)) begin // @[preDebug.scala 25:43]
          bjp_5 <= _GEN_29;
        end
      end
    end
    if (reset) begin // @[preDebug.scala 17:20]
      bjp_6 <= 32'h0; // @[preDebug.scala 17:20]
    end else if (io_IFDone & io_memDone) begin // @[preDebug.scala 19:31]
      if (!(io_exeBranch == 3'h1)) begin // @[preDebug.scala 20:36]
        if (io_exeBranch == 3'h2) begin // @[preDebug.scala 25:43]
          bjp_6 <= _GEN_3;
        end
      end
    end
    if (reset) begin // @[preDebug.scala 18:24]
      bjpMiss_0 <= 32'h0; // @[preDebug.scala 18:24]
    end else if (io_IFDone & io_memDone) begin // @[preDebug.scala 19:31]
      if (io_exeBranch == 3'h1) begin // @[preDebug.scala 20:36]
        if (io_takenMiss) begin // @[preDebug.scala 22:24]
          bjpMiss_0 <= _bjpMiss_0_T_1; // @[preDebug.scala 23:18]
        end
      end
    end
    if (reset) begin // @[preDebug.scala 18:24]
      bjpMiss_1 <= 32'h0; // @[preDebug.scala 18:24]
    end else if (io_IFDone & io_memDone) begin // @[preDebug.scala 19:31]
      if (!(io_exeBranch == 3'h1)) begin // @[preDebug.scala 20:36]
        if (io_exeBranch == 3'h2) begin // @[preDebug.scala 25:43]
          bjpMiss_1 <= _GEN_6;
        end
      end
    end
    if (reset) begin // @[preDebug.scala 18:24]
      bjpMiss_2 <= 32'h0; // @[preDebug.scala 18:24]
    end else if (io_IFDone & io_memDone) begin // @[preDebug.scala 19:31]
      if (!(io_exeBranch == 3'h1)) begin // @[preDebug.scala 20:36]
        if (!(io_exeBranch == 3'h2)) begin // @[preDebug.scala 25:43]
          bjpMiss_2 <= _GEN_24;
        end
      end
    end
    if (reset) begin // @[preDebug.scala 18:24]
      bjpMiss_3 <= 32'h0; // @[preDebug.scala 18:24]
    end else if (io_IFDone & io_memDone) begin // @[preDebug.scala 19:31]
      if (!(io_exeBranch == 3'h1)) begin // @[preDebug.scala 20:36]
        if (!(io_exeBranch == 3'h2)) begin // @[preDebug.scala 25:43]
          bjpMiss_3 <= _GEN_26;
        end
      end
    end
    if (reset) begin // @[preDebug.scala 18:24]
      bjpMiss_4 <= 32'h0; // @[preDebug.scala 18:24]
    end else if (io_IFDone & io_memDone) begin // @[preDebug.scala 19:31]
      if (!(io_exeBranch == 3'h1)) begin // @[preDebug.scala 20:36]
        if (!(io_exeBranch == 3'h2)) begin // @[preDebug.scala 25:43]
          bjpMiss_4 <= _GEN_28;
        end
      end
    end
    if (reset) begin // @[preDebug.scala 18:24]
      bjpMiss_5 <= 32'h0; // @[preDebug.scala 18:24]
    end else if (io_IFDone & io_memDone) begin // @[preDebug.scala 19:31]
      if (!(io_exeBranch == 3'h1)) begin // @[preDebug.scala 20:36]
        if (!(io_exeBranch == 3'h2)) begin // @[preDebug.scala 25:43]
          bjpMiss_5 <= _GEN_30;
        end
      end
    end
    if (reset) begin // @[preDebug.scala 18:24]
      bjpMiss_6 <= 32'h0; // @[preDebug.scala 18:24]
    end else if (io_IFDone & io_memDone) begin // @[preDebug.scala 19:31]
      if (!(io_exeBranch == 3'h1)) begin // @[preDebug.scala 20:36]
        if (io_exeBranch == 3'h2) begin // @[preDebug.scala 25:43]
          bjpMiss_6 <= _GEN_4;
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_9 & ~reset) begin
          $fwrite(32'h80000002,"Name:\tjal\t\tjalr\t\tret\t\tbeq\t\tbne\t\tblt\t\tbge\n"); // @[preDebug.scala 68:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_9 & _T_11) begin
          $fwrite(32'h80000002,"ALL:\t%d\t%d\t%d\t%d\t%d\t%d\t%d\n",bjp_0,bjp_1,bjp_6,bjp_2,bjp_3,bjp_4,bjp_5); // @[preDebug.scala 69:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_9 & _T_11) begin
          $fwrite(32'h80000002,"Miss:\t%d\t%d\t%d\t%d\t%d\t%d\t%d\n",bjpMiss_0,bjpMiss_1,bjpMiss_6,bjpMiss_2,bjpMiss_3,
            bjpMiss_4,bjpMiss_5); // @[preDebug.scala 70:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  bjp_0 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  bjp_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  bjp_2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  bjp_3 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  bjp_4 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  bjp_5 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  bjp_6 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  bjpMiss_0 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  bjpMiss_1 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  bjpMiss_2 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  bjpMiss_3 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  bjpMiss_4 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  bjpMiss_5 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  bjpMiss_6 = _RAND_13[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Core(
  input          clock,
  input          reset,
  output         io_imem_inst_valid,
  input          io_imem_inst_ready,
  output [31:0]  io_imem_inst_addr,
  input  [31:0]  io_imem_inst_read,
  output         io_dmem_data_valid,
  input          io_dmem_data_ready,
  output         io_dmem_data_req,
  output [31:0]  io_dmem_data_addr,
  output [1:0]   io_dmem_data_size,
  output [7:0]   io_dmem_data_strb,
  input  [63:0]  io_dmem_data_read,
  output [127:0] io_dmem_data_write
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  wire  IF_clock; // @[Core.scala 16:18]
  wire  IF_reset; // @[Core.scala 16:18]
  wire  IF_io_imem_inst_valid; // @[Core.scala 16:18]
  wire  IF_io_imem_inst_ready; // @[Core.scala 16:18]
  wire [31:0] IF_io_imem_inst_addr; // @[Core.scala 16:18]
  wire [31:0] IF_io_imem_inst_read; // @[Core.scala 16:18]
  wire  IF_io_takenValid; // @[Core.scala 16:18]
  wire  IF_io_takenValidJalr; // @[Core.scala 16:18]
  wire  IF_io_takenMiss; // @[Core.scala 16:18]
  wire  IF_io_exTakenPre; // @[Core.scala 16:18]
  wire [31:0] IF_io_takenPC; // @[Core.scala 16:18]
  wire [31:0] IF_io_nextPC; // @[Core.scala 16:18]
  wire  IF_io_stall; // @[Core.scala 16:18]
  wire  IF_io_exc; // @[Core.scala 16:18]
  wire  IF_io_intr; // @[Core.scala 16:18]
  wire  IF_io_out_valid; // @[Core.scala 16:18]
  wire [31:0] IF_io_out_pc; // @[Core.scala 16:18]
  wire [31:0] IF_io_out_inst; // @[Core.scala 16:18]
  wire  IF_io_out_takenPre; // @[Core.scala 16:18]
  wire [31:0] IF_io_out_takenPrePC; // @[Core.scala 16:18]
  wire  IF_io_IFDone; // @[Core.scala 16:18]
  wire  IF_io_preRs1En; // @[Core.scala 16:18]
  wire [4:0] IF_io_preRs1Addr; // @[Core.scala 16:18]
  wire [63:0] IF_io_preRs1Data; // @[Core.scala 16:18]
  wire [63:0] IF_io_preRs1x1Data; // @[Core.scala 16:18]
  wire  IF_io_exeX1En; // @[Core.scala 16:18]
  wire [63:0] IF_io_exeAluRes; // @[Core.scala 16:18]
  wire  IF_io_memX1En; // @[Core.scala 16:18]
  wire [63:0] IF_io_memAluRes; // @[Core.scala 16:18]
  wire  IF_io_wbRdEn; // @[Core.scala 16:18]
  wire [4:0] IF_io_wbRdAddr; // @[Core.scala 16:18]
  wire [63:0] IF_io_wbRdData; // @[Core.scala 16:18]
  wire  IfRegId_clock; // @[Core.scala 17:23]
  wire  IfRegId_reset; // @[Core.scala 17:23]
  wire  IfRegId_io_in_valid; // @[Core.scala 17:23]
  wire [31:0] IfRegId_io_in_pc; // @[Core.scala 17:23]
  wire [31:0] IfRegId_io_in_inst; // @[Core.scala 17:23]
  wire  IfRegId_io_in_typeL; // @[Core.scala 17:23]
  wire  IfRegId_io_in_aluA; // @[Core.scala 17:23]
  wire [1:0] IfRegId_io_in_aluB; // @[Core.scala 17:23]
  wire [3:0] IfRegId_io_in_aluOp; // @[Core.scala 17:23]
  wire [2:0] IfRegId_io_in_branch; // @[Core.scala 17:23]
  wire [1:0] IfRegId_io_in_memtoReg; // @[Core.scala 17:23]
  wire  IfRegId_io_in_memWr; // @[Core.scala 17:23]
  wire [2:0] IfRegId_io_in_memOp; // @[Core.scala 17:23]
  wire [31:0] IfRegId_io_in_memAddr; // @[Core.scala 17:23]
  wire  IfRegId_io_in_rdEn; // @[Core.scala 17:23]
  wire [4:0] IfRegId_io_in_rdAddr; // @[Core.scala 17:23]
  wire [63:0] IfRegId_io_in_rs1Data; // @[Core.scala 17:23]
  wire [63:0] IfRegId_io_in_rs2Data; // @[Core.scala 17:23]
  wire [63:0] IfRegId_io_in_imm; // @[Core.scala 17:23]
  wire [63:0] IfRegId_io_in_aluRes; // @[Core.scala 17:23]
  wire [63:0] IfRegId_io_in_memData; // @[Core.scala 17:23]
  wire [3:0] IfRegId_io_in_csrOp; // @[Core.scala 17:23]
  wire  IfRegId_io_in_takenPre; // @[Core.scala 17:23]
  wire [31:0] IfRegId_io_in_takenPrePC; // @[Core.scala 17:23]
  wire  IfRegId_io_out_valid; // @[Core.scala 17:23]
  wire [31:0] IfRegId_io_out_pc; // @[Core.scala 17:23]
  wire [31:0] IfRegId_io_out_inst; // @[Core.scala 17:23]
  wire  IfRegId_io_out_typeL; // @[Core.scala 17:23]
  wire  IfRegId_io_out_aluA; // @[Core.scala 17:23]
  wire [1:0] IfRegId_io_out_aluB; // @[Core.scala 17:23]
  wire [3:0] IfRegId_io_out_aluOp; // @[Core.scala 17:23]
  wire [2:0] IfRegId_io_out_branch; // @[Core.scala 17:23]
  wire [1:0] IfRegId_io_out_memtoReg; // @[Core.scala 17:23]
  wire  IfRegId_io_out_memWr; // @[Core.scala 17:23]
  wire [2:0] IfRegId_io_out_memOp; // @[Core.scala 17:23]
  wire [31:0] IfRegId_io_out_memAddr; // @[Core.scala 17:23]
  wire  IfRegId_io_out_rdEn; // @[Core.scala 17:23]
  wire [4:0] IfRegId_io_out_rdAddr; // @[Core.scala 17:23]
  wire [63:0] IfRegId_io_out_rs1Data; // @[Core.scala 17:23]
  wire [63:0] IfRegId_io_out_rs2Data; // @[Core.scala 17:23]
  wire [63:0] IfRegId_io_out_imm; // @[Core.scala 17:23]
  wire [63:0] IfRegId_io_out_aluRes; // @[Core.scala 17:23]
  wire [63:0] IfRegId_io_out_memData; // @[Core.scala 17:23]
  wire [3:0] IfRegId_io_out_csrOp; // @[Core.scala 17:23]
  wire  IfRegId_io_out_takenPre; // @[Core.scala 17:23]
  wire [31:0] IfRegId_io_out_takenPrePC; // @[Core.scala 17:23]
  wire  IfRegId_io_flush; // @[Core.scala 17:23]
  wire  IfRegId_io_stall; // @[Core.scala 17:23]
  wire  ID_clock; // @[Core.scala 18:18]
  wire  ID_reset; // @[Core.scala 18:18]
  wire  ID_io_rdEn; // @[Core.scala 18:18]
  wire [4:0] ID_io_rdAddr; // @[Core.scala 18:18]
  wire [63:0] ID_io_rdData; // @[Core.scala 18:18]
  wire  ID_io_preRs1En; // @[Core.scala 18:18]
  wire [4:0] ID_io_preRs1Addr; // @[Core.scala 18:18]
  wire [63:0] ID_io_preRs1Data; // @[Core.scala 18:18]
  wire [63:0] ID_io_preRs1x1Data; // @[Core.scala 18:18]
  wire  ID_io_in_valid; // @[Core.scala 18:18]
  wire [31:0] ID_io_in_pc; // @[Core.scala 18:18]
  wire [31:0] ID_io_in_inst; // @[Core.scala 18:18]
  wire  ID_io_in_takenPre; // @[Core.scala 18:18]
  wire [31:0] ID_io_in_takenPrePC; // @[Core.scala 18:18]
  wire  ID_io_exeRdEn; // @[Core.scala 18:18]
  wire [4:0] ID_io_exeRdAddr; // @[Core.scala 18:18]
  wire [63:0] ID_io_exeRdData; // @[Core.scala 18:18]
  wire  ID_io_memRdEn; // @[Core.scala 18:18]
  wire [4:0] ID_io_memRdAddr; // @[Core.scala 18:18]
  wire [63:0] ID_io_memRdData; // @[Core.scala 18:18]
  wire  ID_io_wbRdEn; // @[Core.scala 18:18]
  wire [4:0] ID_io_wbRdAddr; // @[Core.scala 18:18]
  wire [63:0] ID_io_wbRdData; // @[Core.scala 18:18]
  wire  ID_io_bubbleId; // @[Core.scala 18:18]
  wire  ID_io_sBubbleEx; // @[Core.scala 18:18]
  wire  ID_io_sBubbleMem; // @[Core.scala 18:18]
  wire  ID_io_out_valid; // @[Core.scala 18:18]
  wire [31:0] ID_io_out_pc; // @[Core.scala 18:18]
  wire [31:0] ID_io_out_inst; // @[Core.scala 18:18]
  wire  ID_io_out_typeL; // @[Core.scala 18:18]
  wire  ID_io_out_aluA; // @[Core.scala 18:18]
  wire [1:0] ID_io_out_aluB; // @[Core.scala 18:18]
  wire [3:0] ID_io_out_aluOp; // @[Core.scala 18:18]
  wire [2:0] ID_io_out_branch; // @[Core.scala 18:18]
  wire [1:0] ID_io_out_memtoReg; // @[Core.scala 18:18]
  wire  ID_io_out_memWr; // @[Core.scala 18:18]
  wire [2:0] ID_io_out_memOp; // @[Core.scala 18:18]
  wire  ID_io_out_rdEn; // @[Core.scala 18:18]
  wire [4:0] ID_io_out_rdAddr; // @[Core.scala 18:18]
  wire [63:0] ID_io_out_rs1Data; // @[Core.scala 18:18]
  wire [63:0] ID_io_out_rs2Data; // @[Core.scala 18:18]
  wire [63:0] ID_io_out_imm; // @[Core.scala 18:18]
  wire [3:0] ID_io_out_csrOp; // @[Core.scala 18:18]
  wire  ID_io_out_takenPre; // @[Core.scala 18:18]
  wire [31:0] ID_io_out_takenPrePC; // @[Core.scala 18:18]
  wire [63:0] ID_rf_10; // @[Core.scala 18:18]
  wire  IdRegEx_clock; // @[Core.scala 19:23]
  wire  IdRegEx_reset; // @[Core.scala 19:23]
  wire  IdRegEx_io_in_valid; // @[Core.scala 19:23]
  wire [31:0] IdRegEx_io_in_pc; // @[Core.scala 19:23]
  wire [31:0] IdRegEx_io_in_inst; // @[Core.scala 19:23]
  wire  IdRegEx_io_in_typeL; // @[Core.scala 19:23]
  wire  IdRegEx_io_in_aluA; // @[Core.scala 19:23]
  wire [1:0] IdRegEx_io_in_aluB; // @[Core.scala 19:23]
  wire [3:0] IdRegEx_io_in_aluOp; // @[Core.scala 19:23]
  wire [2:0] IdRegEx_io_in_branch; // @[Core.scala 19:23]
  wire [1:0] IdRegEx_io_in_memtoReg; // @[Core.scala 19:23]
  wire  IdRegEx_io_in_memWr; // @[Core.scala 19:23]
  wire [2:0] IdRegEx_io_in_memOp; // @[Core.scala 19:23]
  wire [31:0] IdRegEx_io_in_memAddr; // @[Core.scala 19:23]
  wire  IdRegEx_io_in_rdEn; // @[Core.scala 19:23]
  wire [4:0] IdRegEx_io_in_rdAddr; // @[Core.scala 19:23]
  wire [63:0] IdRegEx_io_in_rs1Data; // @[Core.scala 19:23]
  wire [63:0] IdRegEx_io_in_rs2Data; // @[Core.scala 19:23]
  wire [63:0] IdRegEx_io_in_imm; // @[Core.scala 19:23]
  wire [63:0] IdRegEx_io_in_aluRes; // @[Core.scala 19:23]
  wire [63:0] IdRegEx_io_in_memData; // @[Core.scala 19:23]
  wire [3:0] IdRegEx_io_in_csrOp; // @[Core.scala 19:23]
  wire  IdRegEx_io_in_takenPre; // @[Core.scala 19:23]
  wire [31:0] IdRegEx_io_in_takenPrePC; // @[Core.scala 19:23]
  wire  IdRegEx_io_out_valid; // @[Core.scala 19:23]
  wire [31:0] IdRegEx_io_out_pc; // @[Core.scala 19:23]
  wire [31:0] IdRegEx_io_out_inst; // @[Core.scala 19:23]
  wire  IdRegEx_io_out_typeL; // @[Core.scala 19:23]
  wire  IdRegEx_io_out_aluA; // @[Core.scala 19:23]
  wire [1:0] IdRegEx_io_out_aluB; // @[Core.scala 19:23]
  wire [3:0] IdRegEx_io_out_aluOp; // @[Core.scala 19:23]
  wire [2:0] IdRegEx_io_out_branch; // @[Core.scala 19:23]
  wire [1:0] IdRegEx_io_out_memtoReg; // @[Core.scala 19:23]
  wire  IdRegEx_io_out_memWr; // @[Core.scala 19:23]
  wire [2:0] IdRegEx_io_out_memOp; // @[Core.scala 19:23]
  wire [31:0] IdRegEx_io_out_memAddr; // @[Core.scala 19:23]
  wire  IdRegEx_io_out_rdEn; // @[Core.scala 19:23]
  wire [4:0] IdRegEx_io_out_rdAddr; // @[Core.scala 19:23]
  wire [63:0] IdRegEx_io_out_rs1Data; // @[Core.scala 19:23]
  wire [63:0] IdRegEx_io_out_rs2Data; // @[Core.scala 19:23]
  wire [63:0] IdRegEx_io_out_imm; // @[Core.scala 19:23]
  wire [63:0] IdRegEx_io_out_aluRes; // @[Core.scala 19:23]
  wire [63:0] IdRegEx_io_out_memData; // @[Core.scala 19:23]
  wire [3:0] IdRegEx_io_out_csrOp; // @[Core.scala 19:23]
  wire  IdRegEx_io_out_takenPre; // @[Core.scala 19:23]
  wire [31:0] IdRegEx_io_out_takenPrePC; // @[Core.scala 19:23]
  wire  IdRegEx_io_flush; // @[Core.scala 19:23]
  wire  IdRegEx_io_stall; // @[Core.scala 19:23]
  wire  EX_io_in_valid; // @[Core.scala 20:18]
  wire [31:0] EX_io_in_pc; // @[Core.scala 20:18]
  wire [31:0] EX_io_in_inst; // @[Core.scala 20:18]
  wire  EX_io_in_typeL; // @[Core.scala 20:18]
  wire  EX_io_in_aluA; // @[Core.scala 20:18]
  wire [1:0] EX_io_in_aluB; // @[Core.scala 20:18]
  wire [3:0] EX_io_in_aluOp; // @[Core.scala 20:18]
  wire [2:0] EX_io_in_branch; // @[Core.scala 20:18]
  wire [1:0] EX_io_in_memtoReg; // @[Core.scala 20:18]
  wire  EX_io_in_memWr; // @[Core.scala 20:18]
  wire [2:0] EX_io_in_memOp; // @[Core.scala 20:18]
  wire  EX_io_in_rdEn; // @[Core.scala 20:18]
  wire [4:0] EX_io_in_rdAddr; // @[Core.scala 20:18]
  wire [63:0] EX_io_in_rs1Data; // @[Core.scala 20:18]
  wire [63:0] EX_io_in_rs2Data; // @[Core.scala 20:18]
  wire [63:0] EX_io_in_imm; // @[Core.scala 20:18]
  wire [3:0] EX_io_in_csrOp; // @[Core.scala 20:18]
  wire  EX_io_in_takenPre; // @[Core.scala 20:18]
  wire [31:0] EX_io_in_takenPrePC; // @[Core.scala 20:18]
  wire  EX_io_out_valid; // @[Core.scala 20:18]
  wire [31:0] EX_io_out_pc; // @[Core.scala 20:18]
  wire [31:0] EX_io_out_inst; // @[Core.scala 20:18]
  wire  EX_io_out_typeL; // @[Core.scala 20:18]
  wire  EX_io_out_aluA; // @[Core.scala 20:18]
  wire [1:0] EX_io_out_aluB; // @[Core.scala 20:18]
  wire [3:0] EX_io_out_aluOp; // @[Core.scala 20:18]
  wire [2:0] EX_io_out_branch; // @[Core.scala 20:18]
  wire [1:0] EX_io_out_memtoReg; // @[Core.scala 20:18]
  wire  EX_io_out_memWr; // @[Core.scala 20:18]
  wire [2:0] EX_io_out_memOp; // @[Core.scala 20:18]
  wire  EX_io_out_rdEn; // @[Core.scala 20:18]
  wire [4:0] EX_io_out_rdAddr; // @[Core.scala 20:18]
  wire [63:0] EX_io_out_rs1Data; // @[Core.scala 20:18]
  wire [63:0] EX_io_out_rs2Data; // @[Core.scala 20:18]
  wire [63:0] EX_io_out_imm; // @[Core.scala 20:18]
  wire [31:0] EX_io_out_nextPC; // @[Core.scala 20:18]
  wire [63:0] EX_io_out_aluRes; // @[Core.scala 20:18]
  wire [3:0] EX_io_out_csrOp; // @[Core.scala 20:18]
  wire  EX_io_out_takenPre; // @[Core.scala 20:18]
  wire [31:0] EX_io_out_takenPrePC; // @[Core.scala 20:18]
  wire [63:0] EX_io_exeRdData; // @[Core.scala 20:18]
  wire  EX_io_bubbleEx; // @[Core.scala 20:18]
  wire  EX_io_takenValid; // @[Core.scala 20:18]
  wire  EX_io_takenValidJalr; // @[Core.scala 20:18]
  wire  EX_io_takenMiss; // @[Core.scala 20:18]
  wire  EX_io_exTakenPre; // @[Core.scala 20:18]
  wire [31:0] EX_io_takenPC; // @[Core.scala 20:18]
  wire  EX_io_exeX1En; // @[Core.scala 20:18]
  wire [63:0] EX_io_exeAluRes; // @[Core.scala 20:18]
  wire  EX_io_exc; // @[Core.scala 20:18]
  wire [3:0] EX_io_csrOp; // @[Core.scala 20:18]
  wire [63:0] EX_io_mepc; // @[Core.scala 20:18]
  wire [63:0] EX_io_mtvec; // @[Core.scala 20:18]
  wire  EX_io_time_int; // @[Core.scala 20:18]
  wire  ExRegMem_clock; // @[Core.scala 21:24]
  wire  ExRegMem_reset; // @[Core.scala 21:24]
  wire  ExRegMem_io_in_valid; // @[Core.scala 21:24]
  wire [31:0] ExRegMem_io_in_pc; // @[Core.scala 21:24]
  wire [31:0] ExRegMem_io_in_inst; // @[Core.scala 21:24]
  wire  ExRegMem_io_in_typeL; // @[Core.scala 21:24]
  wire  ExRegMem_io_in_aluA; // @[Core.scala 21:24]
  wire [1:0] ExRegMem_io_in_aluB; // @[Core.scala 21:24]
  wire [3:0] ExRegMem_io_in_aluOp; // @[Core.scala 21:24]
  wire [2:0] ExRegMem_io_in_branch; // @[Core.scala 21:24]
  wire [1:0] ExRegMem_io_in_memtoReg; // @[Core.scala 21:24]
  wire  ExRegMem_io_in_memWr; // @[Core.scala 21:24]
  wire [2:0] ExRegMem_io_in_memOp; // @[Core.scala 21:24]
  wire [31:0] ExRegMem_io_in_memAddr; // @[Core.scala 21:24]
  wire  ExRegMem_io_in_rdEn; // @[Core.scala 21:24]
  wire [4:0] ExRegMem_io_in_rdAddr; // @[Core.scala 21:24]
  wire [63:0] ExRegMem_io_in_rs1Data; // @[Core.scala 21:24]
  wire [63:0] ExRegMem_io_in_rs2Data; // @[Core.scala 21:24]
  wire [63:0] ExRegMem_io_in_imm; // @[Core.scala 21:24]
  wire [63:0] ExRegMem_io_in_aluRes; // @[Core.scala 21:24]
  wire [63:0] ExRegMem_io_in_memData; // @[Core.scala 21:24]
  wire [3:0] ExRegMem_io_in_csrOp; // @[Core.scala 21:24]
  wire  ExRegMem_io_in_takenPre; // @[Core.scala 21:24]
  wire [31:0] ExRegMem_io_in_takenPrePC; // @[Core.scala 21:24]
  wire  ExRegMem_io_out_valid; // @[Core.scala 21:24]
  wire [31:0] ExRegMem_io_out_pc; // @[Core.scala 21:24]
  wire [31:0] ExRegMem_io_out_inst; // @[Core.scala 21:24]
  wire  ExRegMem_io_out_typeL; // @[Core.scala 21:24]
  wire  ExRegMem_io_out_aluA; // @[Core.scala 21:24]
  wire [1:0] ExRegMem_io_out_aluB; // @[Core.scala 21:24]
  wire [3:0] ExRegMem_io_out_aluOp; // @[Core.scala 21:24]
  wire [2:0] ExRegMem_io_out_branch; // @[Core.scala 21:24]
  wire [1:0] ExRegMem_io_out_memtoReg; // @[Core.scala 21:24]
  wire  ExRegMem_io_out_memWr; // @[Core.scala 21:24]
  wire [2:0] ExRegMem_io_out_memOp; // @[Core.scala 21:24]
  wire [31:0] ExRegMem_io_out_memAddr; // @[Core.scala 21:24]
  wire  ExRegMem_io_out_rdEn; // @[Core.scala 21:24]
  wire [4:0] ExRegMem_io_out_rdAddr; // @[Core.scala 21:24]
  wire [63:0] ExRegMem_io_out_rs1Data; // @[Core.scala 21:24]
  wire [63:0] ExRegMem_io_out_rs2Data; // @[Core.scala 21:24]
  wire [63:0] ExRegMem_io_out_imm; // @[Core.scala 21:24]
  wire [63:0] ExRegMem_io_out_aluRes; // @[Core.scala 21:24]
  wire [63:0] ExRegMem_io_out_memData; // @[Core.scala 21:24]
  wire [3:0] ExRegMem_io_out_csrOp; // @[Core.scala 21:24]
  wire  ExRegMem_io_out_takenPre; // @[Core.scala 21:24]
  wire [31:0] ExRegMem_io_out_takenPrePC; // @[Core.scala 21:24]
  wire  ExRegMem_io_flush; // @[Core.scala 21:24]
  wire  ExRegMem_io_stall; // @[Core.scala 21:24]
  wire  MEM_clock; // @[Core.scala 22:19]
  wire  MEM_reset; // @[Core.scala 22:19]
  wire  MEM_io_dmem_data_valid; // @[Core.scala 22:19]
  wire  MEM_io_dmem_data_ready; // @[Core.scala 22:19]
  wire  MEM_io_dmem_data_req; // @[Core.scala 22:19]
  wire [31:0] MEM_io_dmem_data_addr; // @[Core.scala 22:19]
  wire [1:0] MEM_io_dmem_data_size; // @[Core.scala 22:19]
  wire [7:0] MEM_io_dmem_data_strb; // @[Core.scala 22:19]
  wire [63:0] MEM_io_dmem_data_read; // @[Core.scala 22:19]
  wire [127:0] MEM_io_dmem_data_write; // @[Core.scala 22:19]
  wire  MEM_io_IFDone; // @[Core.scala 22:19]
  wire  MEM_io_in_valid; // @[Core.scala 22:19]
  wire [31:0] MEM_io_in_pc; // @[Core.scala 22:19]
  wire [31:0] MEM_io_in_inst; // @[Core.scala 22:19]
  wire  MEM_io_in_typeL; // @[Core.scala 22:19]
  wire  MEM_io_in_aluA; // @[Core.scala 22:19]
  wire [1:0] MEM_io_in_aluB; // @[Core.scala 22:19]
  wire [3:0] MEM_io_in_aluOp; // @[Core.scala 22:19]
  wire [2:0] MEM_io_in_branch; // @[Core.scala 22:19]
  wire [1:0] MEM_io_in_memtoReg; // @[Core.scala 22:19]
  wire  MEM_io_in_memWr; // @[Core.scala 22:19]
  wire [2:0] MEM_io_in_memOp; // @[Core.scala 22:19]
  wire  MEM_io_in_rdEn; // @[Core.scala 22:19]
  wire [4:0] MEM_io_in_rdAddr; // @[Core.scala 22:19]
  wire [63:0] MEM_io_in_rs1Data; // @[Core.scala 22:19]
  wire [63:0] MEM_io_in_rs2Data; // @[Core.scala 22:19]
  wire [63:0] MEM_io_in_imm; // @[Core.scala 22:19]
  wire [63:0] MEM_io_in_aluRes; // @[Core.scala 22:19]
  wire [3:0] MEM_io_in_csrOp; // @[Core.scala 22:19]
  wire  MEM_io_in_takenPre; // @[Core.scala 22:19]
  wire [31:0] MEM_io_in_takenPrePC; // @[Core.scala 22:19]
  wire  MEM_io_out_valid; // @[Core.scala 22:19]
  wire [31:0] MEM_io_out_pc; // @[Core.scala 22:19]
  wire [31:0] MEM_io_out_inst; // @[Core.scala 22:19]
  wire  MEM_io_out_typeL; // @[Core.scala 22:19]
  wire  MEM_io_out_aluA; // @[Core.scala 22:19]
  wire [1:0] MEM_io_out_aluB; // @[Core.scala 22:19]
  wire [3:0] MEM_io_out_aluOp; // @[Core.scala 22:19]
  wire [2:0] MEM_io_out_branch; // @[Core.scala 22:19]
  wire [1:0] MEM_io_out_memtoReg; // @[Core.scala 22:19]
  wire  MEM_io_out_memWr; // @[Core.scala 22:19]
  wire [2:0] MEM_io_out_memOp; // @[Core.scala 22:19]
  wire [31:0] MEM_io_out_memAddr; // @[Core.scala 22:19]
  wire  MEM_io_out_rdEn; // @[Core.scala 22:19]
  wire [4:0] MEM_io_out_rdAddr; // @[Core.scala 22:19]
  wire [63:0] MEM_io_out_rs1Data; // @[Core.scala 22:19]
  wire [63:0] MEM_io_out_rs2Data; // @[Core.scala 22:19]
  wire [63:0] MEM_io_out_imm; // @[Core.scala 22:19]
  wire [63:0] MEM_io_out_aluRes; // @[Core.scala 22:19]
  wire [63:0] MEM_io_out_memData; // @[Core.scala 22:19]
  wire [3:0] MEM_io_out_csrOp; // @[Core.scala 22:19]
  wire  MEM_io_out_takenPre; // @[Core.scala 22:19]
  wire [31:0] MEM_io_out_takenPrePC; // @[Core.scala 22:19]
  wire [63:0] MEM_io_memRdData; // @[Core.scala 22:19]
  wire  MEM_io_memDone; // @[Core.scala 22:19]
  wire  MEM_io_memX1En; // @[Core.scala 22:19]
  wire [63:0] MEM_io_memAluRes; // @[Core.scala 22:19]
  wire  MEM_io_cmp_ren; // @[Core.scala 22:19]
  wire  MEM_io_cmp_wen; // @[Core.scala 22:19]
  wire [63:0] MEM_io_cmp_addr; // @[Core.scala 22:19]
  wire [63:0] MEM_io_cmp_wdata; // @[Core.scala 22:19]
  wire [63:0] MEM_io_cmp_rdata; // @[Core.scala 22:19]
  wire  MemRegWb_clock; // @[Core.scala 23:24]
  wire  MemRegWb_reset; // @[Core.scala 23:24]
  wire  MemRegWb_io_in_valid; // @[Core.scala 23:24]
  wire [31:0] MemRegWb_io_in_pc; // @[Core.scala 23:24]
  wire [31:0] MemRegWb_io_in_inst; // @[Core.scala 23:24]
  wire  MemRegWb_io_in_typeL; // @[Core.scala 23:24]
  wire  MemRegWb_io_in_aluA; // @[Core.scala 23:24]
  wire [1:0] MemRegWb_io_in_aluB; // @[Core.scala 23:24]
  wire [3:0] MemRegWb_io_in_aluOp; // @[Core.scala 23:24]
  wire [2:0] MemRegWb_io_in_branch; // @[Core.scala 23:24]
  wire [1:0] MemRegWb_io_in_memtoReg; // @[Core.scala 23:24]
  wire  MemRegWb_io_in_memWr; // @[Core.scala 23:24]
  wire [2:0] MemRegWb_io_in_memOp; // @[Core.scala 23:24]
  wire [31:0] MemRegWb_io_in_memAddr; // @[Core.scala 23:24]
  wire  MemRegWb_io_in_rdEn; // @[Core.scala 23:24]
  wire [4:0] MemRegWb_io_in_rdAddr; // @[Core.scala 23:24]
  wire [63:0] MemRegWb_io_in_rs1Data; // @[Core.scala 23:24]
  wire [63:0] MemRegWb_io_in_rs2Data; // @[Core.scala 23:24]
  wire [63:0] MemRegWb_io_in_imm; // @[Core.scala 23:24]
  wire [63:0] MemRegWb_io_in_aluRes; // @[Core.scala 23:24]
  wire [63:0] MemRegWb_io_in_memData; // @[Core.scala 23:24]
  wire [3:0] MemRegWb_io_in_csrOp; // @[Core.scala 23:24]
  wire  MemRegWb_io_in_takenPre; // @[Core.scala 23:24]
  wire [31:0] MemRegWb_io_in_takenPrePC; // @[Core.scala 23:24]
  wire  MemRegWb_io_out_valid; // @[Core.scala 23:24]
  wire [31:0] MemRegWb_io_out_pc; // @[Core.scala 23:24]
  wire [31:0] MemRegWb_io_out_inst; // @[Core.scala 23:24]
  wire  MemRegWb_io_out_typeL; // @[Core.scala 23:24]
  wire  MemRegWb_io_out_aluA; // @[Core.scala 23:24]
  wire [1:0] MemRegWb_io_out_aluB; // @[Core.scala 23:24]
  wire [3:0] MemRegWb_io_out_aluOp; // @[Core.scala 23:24]
  wire [2:0] MemRegWb_io_out_branch; // @[Core.scala 23:24]
  wire [1:0] MemRegWb_io_out_memtoReg; // @[Core.scala 23:24]
  wire  MemRegWb_io_out_memWr; // @[Core.scala 23:24]
  wire [2:0] MemRegWb_io_out_memOp; // @[Core.scala 23:24]
  wire [31:0] MemRegWb_io_out_memAddr; // @[Core.scala 23:24]
  wire  MemRegWb_io_out_rdEn; // @[Core.scala 23:24]
  wire [4:0] MemRegWb_io_out_rdAddr; // @[Core.scala 23:24]
  wire [63:0] MemRegWb_io_out_rs1Data; // @[Core.scala 23:24]
  wire [63:0] MemRegWb_io_out_rs2Data; // @[Core.scala 23:24]
  wire [63:0] MemRegWb_io_out_imm; // @[Core.scala 23:24]
  wire [63:0] MemRegWb_io_out_aluRes; // @[Core.scala 23:24]
  wire [63:0] MemRegWb_io_out_memData; // @[Core.scala 23:24]
  wire [3:0] MemRegWb_io_out_csrOp; // @[Core.scala 23:24]
  wire  MemRegWb_io_out_takenPre; // @[Core.scala 23:24]
  wire [31:0] MemRegWb_io_out_takenPrePC; // @[Core.scala 23:24]
  wire  MemRegWb_io_flush; // @[Core.scala 23:24]
  wire  MemRegWb_io_stall; // @[Core.scala 23:24]
  wire  WB_clock; // @[Core.scala 24:18]
  wire  WB_reset; // @[Core.scala 24:18]
  wire  WB_io_in_valid; // @[Core.scala 24:18]
  wire [31:0] WB_io_in_pc; // @[Core.scala 24:18]
  wire [31:0] WB_io_in_inst; // @[Core.scala 24:18]
  wire [1:0] WB_io_in_memtoReg; // @[Core.scala 24:18]
  wire  WB_io_in_memWr; // @[Core.scala 24:18]
  wire [31:0] WB_io_in_memAddr; // @[Core.scala 24:18]
  wire  WB_io_in_rdEn; // @[Core.scala 24:18]
  wire [4:0] WB_io_in_rdAddr; // @[Core.scala 24:18]
  wire [63:0] WB_io_in_rs1Data; // @[Core.scala 24:18]
  wire [63:0] WB_io_in_aluRes; // @[Core.scala 24:18]
  wire [63:0] WB_io_in_memData; // @[Core.scala 24:18]
  wire [3:0] WB_io_in_csrOp; // @[Core.scala 24:18]
  wire  WB_io_IFDone; // @[Core.scala 24:18]
  wire  WB_io_memDone; // @[Core.scala 24:18]
  wire [31:0] WB_io_pc_intr; // @[Core.scala 24:18]
  wire [31:0] WB_io_pc; // @[Core.scala 24:18]
  wire [31:0] WB_io_inst; // @[Core.scala 24:18]
  wire  WB_io_wbRdEn; // @[Core.scala 24:18]
  wire [4:0] WB_io_wbRdAddr; // @[Core.scala 24:18]
  wire [63:0] WB_io_wbRdData; // @[Core.scala 24:18]
  wire  WB_io_ready_cmt; // @[Core.scala 24:18]
  wire [3:0] WB_io_csrOp_WB; // @[Core.scala 24:18]
  wire [63:0] WB_io_mepc; // @[Core.scala 24:18]
  wire [63:0] WB_io_mtvec; // @[Core.scala 24:18]
  wire  WB_io_cmp_ren; // @[Core.scala 24:18]
  wire  WB_io_cmp_wen; // @[Core.scala 24:18]
  wire [63:0] WB_io_cmp_addr; // @[Core.scala 24:18]
  wire [63:0] WB_io_cmp_wdata; // @[Core.scala 24:18]
  wire [63:0] WB_io_cmp_rdata; // @[Core.scala 24:18]
  wire  WB_io_exc; // @[Core.scala 24:18]
  wire [1:0] WB_io_memtoReg; // @[Core.scala 24:18]
  wire  WB_io_memWr; // @[Core.scala 24:18]
  wire [31:0] WB_io_mem_addr; // @[Core.scala 24:18]
  wire  WB_io_time_int; // @[Core.scala 24:18]
  wire  preDebug_clock; // @[Core.scala 27:24]
  wire  preDebug_reset; // @[Core.scala 27:24]
  wire [2:0] preDebug_io_exeBranch; // @[Core.scala 27:24]
  wire  preDebug_io_takenMiss; // @[Core.scala 27:24]
  wire [4:0] preDebug_io_rs1Addr; // @[Core.scala 27:24]
  wire  preDebug_io_coreEnd; // @[Core.scala 27:24]
  wire  preDebug_io_IFDone; // @[Core.scala 27:24]
  wire  preDebug_io_memDone; // @[Core.scala 27:24]
  wire  dt_ic_clock; // @[Core.scala 166:21]
  wire [7:0] dt_ic_coreid; // @[Core.scala 166:21]
  wire [7:0] dt_ic_index; // @[Core.scala 166:21]
  wire  dt_ic_valid; // @[Core.scala 166:21]
  wire [63:0] dt_ic_pc; // @[Core.scala 166:21]
  wire [31:0] dt_ic_instr; // @[Core.scala 166:21]
  wire  dt_ic_skip; // @[Core.scala 166:21]
  wire  dt_ic_isRVC; // @[Core.scala 166:21]
  wire  dt_ic_scFailed; // @[Core.scala 166:21]
  wire  dt_ic_wen; // @[Core.scala 166:21]
  wire [63:0] dt_ic_wdata; // @[Core.scala 166:21]
  wire [7:0] dt_ic_wdest; // @[Core.scala 166:21]
  wire  dt_ae_clock; // @[Core.scala 180:21]
  wire [7:0] dt_ae_coreid; // @[Core.scala 180:21]
  wire [31:0] dt_ae_intrNO; // @[Core.scala 180:21]
  wire [31:0] dt_ae_cause; // @[Core.scala 180:21]
  wire [63:0] dt_ae_exceptionPC; // @[Core.scala 180:21]
  wire [31:0] dt_ae_exceptionInst; // @[Core.scala 180:21]
  wire  dt_te_clock; // @[Core.scala 193:21]
  wire [7:0] dt_te_coreid; // @[Core.scala 193:21]
  wire  dt_te_valid; // @[Core.scala 193:21]
  wire [2:0] dt_te_code; // @[Core.scala 193:21]
  wire [63:0] dt_te_pc; // @[Core.scala 193:21]
  wire [63:0] dt_te_cycleCnt; // @[Core.scala 193:21]
  wire [63:0] dt_te_instrCnt; // @[Core.scala 193:21]
  wire [31:0] _exceptionPC_T_4 = ID_io_out_pc != 32'h0 ? ID_io_out_pc : IF_io_out_pc; // @[Core.scala 40:40]
  wire [31:0] _exceptionPC_T_5 = EX_io_out_pc != 32'h0 ? EX_io_out_pc : _exceptionPC_T_4; // @[Core.scala 39:38]
  wire [31:0] _exceptionPC_T_6 = MEM_io_out_pc != 32'h0 ? MEM_io_out_pc : _exceptionPC_T_5; // @[Core.scala 38:36]
  wire [31:0] _exceptionPC_T_7 = WB_io_pc != 32'h0 ? WB_io_pc : _exceptionPC_T_6; // @[Core.scala 37:34]
  wire  EXLHitID = ID_io_bubbleId & EX_io_bubbleEx; // @[Core.scala 43:33]
  wire  EXSHitID = ID_io_sBubbleEx & EX_io_out_csrOp != 4'h0; // @[Core.scala 46:34]
  wire  MEMSHitID = ID_io_sBubbleMem & MEM_io_out_csrOp != 4'h0; // @[Core.scala 47:36]
  wire  EXSHitIDEn = EXSHitID | MEMSHitID; // @[Core.scala 48:29]
  wire  ecallEn = WB_io_csrOp_WB[3] | WB_io_time_int; // @[Core.scala 50:43]
  wire  _stallIfIdEn_T = ~IF_io_IFDone; // @[Core.scala 59:22]
  wire  _stallIfIdEn_T_1 = ~MEM_io_memDone; // @[Core.scala 59:39]
  wire  valid = WB_io_ready_cmt & IF_io_IFDone & MEM_io_memDone; // @[Core.scala 153:47]
  wire [31:0] _T = WB_io_inst; // @[Core.scala 158:20]
  wire  _T_1 = 32'h7b == _T; // @[Core.scala 158:20]
  wire  _T_2 = 32'h7b == _T & valid; // @[Core.scala 158:32]
  wire  _req_clint_T_5 = WB_io_memtoReg == 2'h1 | WB_io_memWr; // @[Core.scala 163:43]
  wire  req_clint = (WB_io_mem_addr == 32'h2004000 | WB_io_mem_addr == 32'h200bff8) & _req_clint_T_5; // @[Core.scala 162:77]
  reg  dt_ic_io_valid_REG; // @[Core.scala 170:31]
  reg [31:0] dt_ic_io_pc_REG; // @[Core.scala 171:31]
  reg [31:0] dt_ic_io_instr_REG; // @[Core.scala 172:31]
  reg  dt_ic_io_skip_REG; // @[Core.scala 173:31]
  reg  dt_ic_io_wen_REG; // @[Core.scala 176:31]
  reg [63:0] dt_ic_io_wdata_REG; // @[Core.scala 177:31]
  reg [4:0] dt_ic_io_wdest_REG; // @[Core.scala 178:31]
  reg [2:0] dt_ae_io_intrNO_REG; // @[Core.scala 183:35]
  reg [31:0] dt_ae_io_exceptionPC_REG; // @[Core.scala 185:35]
  reg [63:0] cycle_cnt; // @[Core.scala 187:26]
  reg [63:0] instr_cnt; // @[Core.scala 188:26]
  wire [63:0] _cycle_cnt_T_1 = cycle_cnt + 64'h1; // @[Core.scala 190:26]
  wire [63:0] _GEN_0 = {{63'd0}, valid}; // @[Core.scala 191:26]
  wire [63:0] _instr_cnt_T_1 = instr_cnt + _GEN_0; // @[Core.scala 191:26]
  wire [63:0] rf_a0_0 = ID_rf_10;
  InstFetch IF ( // @[Core.scala 16:18]
    .clock(IF_clock),
    .reset(IF_reset),
    .io_imem_inst_valid(IF_io_imem_inst_valid),
    .io_imem_inst_ready(IF_io_imem_inst_ready),
    .io_imem_inst_addr(IF_io_imem_inst_addr),
    .io_imem_inst_read(IF_io_imem_inst_read),
    .io_takenValid(IF_io_takenValid),
    .io_takenValidJalr(IF_io_takenValidJalr),
    .io_takenMiss(IF_io_takenMiss),
    .io_exTakenPre(IF_io_exTakenPre),
    .io_takenPC(IF_io_takenPC),
    .io_nextPC(IF_io_nextPC),
    .io_stall(IF_io_stall),
    .io_exc(IF_io_exc),
    .io_intr(IF_io_intr),
    .io_out_valid(IF_io_out_valid),
    .io_out_pc(IF_io_out_pc),
    .io_out_inst(IF_io_out_inst),
    .io_out_takenPre(IF_io_out_takenPre),
    .io_out_takenPrePC(IF_io_out_takenPrePC),
    .io_IFDone(IF_io_IFDone),
    .io_preRs1En(IF_io_preRs1En),
    .io_preRs1Addr(IF_io_preRs1Addr),
    .io_preRs1Data(IF_io_preRs1Data),
    .io_preRs1x1Data(IF_io_preRs1x1Data),
    .io_exeX1En(IF_io_exeX1En),
    .io_exeAluRes(IF_io_exeAluRes),
    .io_memX1En(IF_io_memX1En),
    .io_memAluRes(IF_io_memAluRes),
    .io_wbRdEn(IF_io_wbRdEn),
    .io_wbRdAddr(IF_io_wbRdAddr),
    .io_wbRdData(IF_io_wbRdData)
  );
  PipelineReg IfRegId ( // @[Core.scala 17:23]
    .clock(IfRegId_clock),
    .reset(IfRegId_reset),
    .io_in_valid(IfRegId_io_in_valid),
    .io_in_pc(IfRegId_io_in_pc),
    .io_in_inst(IfRegId_io_in_inst),
    .io_in_typeL(IfRegId_io_in_typeL),
    .io_in_aluA(IfRegId_io_in_aluA),
    .io_in_aluB(IfRegId_io_in_aluB),
    .io_in_aluOp(IfRegId_io_in_aluOp),
    .io_in_branch(IfRegId_io_in_branch),
    .io_in_memtoReg(IfRegId_io_in_memtoReg),
    .io_in_memWr(IfRegId_io_in_memWr),
    .io_in_memOp(IfRegId_io_in_memOp),
    .io_in_memAddr(IfRegId_io_in_memAddr),
    .io_in_rdEn(IfRegId_io_in_rdEn),
    .io_in_rdAddr(IfRegId_io_in_rdAddr),
    .io_in_rs1Data(IfRegId_io_in_rs1Data),
    .io_in_rs2Data(IfRegId_io_in_rs2Data),
    .io_in_imm(IfRegId_io_in_imm),
    .io_in_aluRes(IfRegId_io_in_aluRes),
    .io_in_memData(IfRegId_io_in_memData),
    .io_in_csrOp(IfRegId_io_in_csrOp),
    .io_in_takenPre(IfRegId_io_in_takenPre),
    .io_in_takenPrePC(IfRegId_io_in_takenPrePC),
    .io_out_valid(IfRegId_io_out_valid),
    .io_out_pc(IfRegId_io_out_pc),
    .io_out_inst(IfRegId_io_out_inst),
    .io_out_typeL(IfRegId_io_out_typeL),
    .io_out_aluA(IfRegId_io_out_aluA),
    .io_out_aluB(IfRegId_io_out_aluB),
    .io_out_aluOp(IfRegId_io_out_aluOp),
    .io_out_branch(IfRegId_io_out_branch),
    .io_out_memtoReg(IfRegId_io_out_memtoReg),
    .io_out_memWr(IfRegId_io_out_memWr),
    .io_out_memOp(IfRegId_io_out_memOp),
    .io_out_memAddr(IfRegId_io_out_memAddr),
    .io_out_rdEn(IfRegId_io_out_rdEn),
    .io_out_rdAddr(IfRegId_io_out_rdAddr),
    .io_out_rs1Data(IfRegId_io_out_rs1Data),
    .io_out_rs2Data(IfRegId_io_out_rs2Data),
    .io_out_imm(IfRegId_io_out_imm),
    .io_out_aluRes(IfRegId_io_out_aluRes),
    .io_out_memData(IfRegId_io_out_memData),
    .io_out_csrOp(IfRegId_io_out_csrOp),
    .io_out_takenPre(IfRegId_io_out_takenPre),
    .io_out_takenPrePC(IfRegId_io_out_takenPrePC),
    .io_flush(IfRegId_io_flush),
    .io_stall(IfRegId_io_stall)
  );
  Decode ID ( // @[Core.scala 18:18]
    .clock(ID_clock),
    .reset(ID_reset),
    .io_rdEn(ID_io_rdEn),
    .io_rdAddr(ID_io_rdAddr),
    .io_rdData(ID_io_rdData),
    .io_preRs1En(ID_io_preRs1En),
    .io_preRs1Addr(ID_io_preRs1Addr),
    .io_preRs1Data(ID_io_preRs1Data),
    .io_preRs1x1Data(ID_io_preRs1x1Data),
    .io_in_valid(ID_io_in_valid),
    .io_in_pc(ID_io_in_pc),
    .io_in_inst(ID_io_in_inst),
    .io_in_takenPre(ID_io_in_takenPre),
    .io_in_takenPrePC(ID_io_in_takenPrePC),
    .io_exeRdEn(ID_io_exeRdEn),
    .io_exeRdAddr(ID_io_exeRdAddr),
    .io_exeRdData(ID_io_exeRdData),
    .io_memRdEn(ID_io_memRdEn),
    .io_memRdAddr(ID_io_memRdAddr),
    .io_memRdData(ID_io_memRdData),
    .io_wbRdEn(ID_io_wbRdEn),
    .io_wbRdAddr(ID_io_wbRdAddr),
    .io_wbRdData(ID_io_wbRdData),
    .io_bubbleId(ID_io_bubbleId),
    .io_sBubbleEx(ID_io_sBubbleEx),
    .io_sBubbleMem(ID_io_sBubbleMem),
    .io_out_valid(ID_io_out_valid),
    .io_out_pc(ID_io_out_pc),
    .io_out_inst(ID_io_out_inst),
    .io_out_typeL(ID_io_out_typeL),
    .io_out_aluA(ID_io_out_aluA),
    .io_out_aluB(ID_io_out_aluB),
    .io_out_aluOp(ID_io_out_aluOp),
    .io_out_branch(ID_io_out_branch),
    .io_out_memtoReg(ID_io_out_memtoReg),
    .io_out_memWr(ID_io_out_memWr),
    .io_out_memOp(ID_io_out_memOp),
    .io_out_rdEn(ID_io_out_rdEn),
    .io_out_rdAddr(ID_io_out_rdAddr),
    .io_out_rs1Data(ID_io_out_rs1Data),
    .io_out_rs2Data(ID_io_out_rs2Data),
    .io_out_imm(ID_io_out_imm),
    .io_out_csrOp(ID_io_out_csrOp),
    .io_out_takenPre(ID_io_out_takenPre),
    .io_out_takenPrePC(ID_io_out_takenPrePC),
    .rf_10(ID_rf_10)
  );
  PipelineReg IdRegEx ( // @[Core.scala 19:23]
    .clock(IdRegEx_clock),
    .reset(IdRegEx_reset),
    .io_in_valid(IdRegEx_io_in_valid),
    .io_in_pc(IdRegEx_io_in_pc),
    .io_in_inst(IdRegEx_io_in_inst),
    .io_in_typeL(IdRegEx_io_in_typeL),
    .io_in_aluA(IdRegEx_io_in_aluA),
    .io_in_aluB(IdRegEx_io_in_aluB),
    .io_in_aluOp(IdRegEx_io_in_aluOp),
    .io_in_branch(IdRegEx_io_in_branch),
    .io_in_memtoReg(IdRegEx_io_in_memtoReg),
    .io_in_memWr(IdRegEx_io_in_memWr),
    .io_in_memOp(IdRegEx_io_in_memOp),
    .io_in_memAddr(IdRegEx_io_in_memAddr),
    .io_in_rdEn(IdRegEx_io_in_rdEn),
    .io_in_rdAddr(IdRegEx_io_in_rdAddr),
    .io_in_rs1Data(IdRegEx_io_in_rs1Data),
    .io_in_rs2Data(IdRegEx_io_in_rs2Data),
    .io_in_imm(IdRegEx_io_in_imm),
    .io_in_aluRes(IdRegEx_io_in_aluRes),
    .io_in_memData(IdRegEx_io_in_memData),
    .io_in_csrOp(IdRegEx_io_in_csrOp),
    .io_in_takenPre(IdRegEx_io_in_takenPre),
    .io_in_takenPrePC(IdRegEx_io_in_takenPrePC),
    .io_out_valid(IdRegEx_io_out_valid),
    .io_out_pc(IdRegEx_io_out_pc),
    .io_out_inst(IdRegEx_io_out_inst),
    .io_out_typeL(IdRegEx_io_out_typeL),
    .io_out_aluA(IdRegEx_io_out_aluA),
    .io_out_aluB(IdRegEx_io_out_aluB),
    .io_out_aluOp(IdRegEx_io_out_aluOp),
    .io_out_branch(IdRegEx_io_out_branch),
    .io_out_memtoReg(IdRegEx_io_out_memtoReg),
    .io_out_memWr(IdRegEx_io_out_memWr),
    .io_out_memOp(IdRegEx_io_out_memOp),
    .io_out_memAddr(IdRegEx_io_out_memAddr),
    .io_out_rdEn(IdRegEx_io_out_rdEn),
    .io_out_rdAddr(IdRegEx_io_out_rdAddr),
    .io_out_rs1Data(IdRegEx_io_out_rs1Data),
    .io_out_rs2Data(IdRegEx_io_out_rs2Data),
    .io_out_imm(IdRegEx_io_out_imm),
    .io_out_aluRes(IdRegEx_io_out_aluRes),
    .io_out_memData(IdRegEx_io_out_memData),
    .io_out_csrOp(IdRegEx_io_out_csrOp),
    .io_out_takenPre(IdRegEx_io_out_takenPre),
    .io_out_takenPrePC(IdRegEx_io_out_takenPrePC),
    .io_flush(IdRegEx_io_flush),
    .io_stall(IdRegEx_io_stall)
  );
  Execution EX ( // @[Core.scala 20:18]
    .io_in_valid(EX_io_in_valid),
    .io_in_pc(EX_io_in_pc),
    .io_in_inst(EX_io_in_inst),
    .io_in_typeL(EX_io_in_typeL),
    .io_in_aluA(EX_io_in_aluA),
    .io_in_aluB(EX_io_in_aluB),
    .io_in_aluOp(EX_io_in_aluOp),
    .io_in_branch(EX_io_in_branch),
    .io_in_memtoReg(EX_io_in_memtoReg),
    .io_in_memWr(EX_io_in_memWr),
    .io_in_memOp(EX_io_in_memOp),
    .io_in_rdEn(EX_io_in_rdEn),
    .io_in_rdAddr(EX_io_in_rdAddr),
    .io_in_rs1Data(EX_io_in_rs1Data),
    .io_in_rs2Data(EX_io_in_rs2Data),
    .io_in_imm(EX_io_in_imm),
    .io_in_csrOp(EX_io_in_csrOp),
    .io_in_takenPre(EX_io_in_takenPre),
    .io_in_takenPrePC(EX_io_in_takenPrePC),
    .io_out_valid(EX_io_out_valid),
    .io_out_pc(EX_io_out_pc),
    .io_out_inst(EX_io_out_inst),
    .io_out_typeL(EX_io_out_typeL),
    .io_out_aluA(EX_io_out_aluA),
    .io_out_aluB(EX_io_out_aluB),
    .io_out_aluOp(EX_io_out_aluOp),
    .io_out_branch(EX_io_out_branch),
    .io_out_memtoReg(EX_io_out_memtoReg),
    .io_out_memWr(EX_io_out_memWr),
    .io_out_memOp(EX_io_out_memOp),
    .io_out_rdEn(EX_io_out_rdEn),
    .io_out_rdAddr(EX_io_out_rdAddr),
    .io_out_rs1Data(EX_io_out_rs1Data),
    .io_out_rs2Data(EX_io_out_rs2Data),
    .io_out_imm(EX_io_out_imm),
    .io_out_nextPC(EX_io_out_nextPC),
    .io_out_aluRes(EX_io_out_aluRes),
    .io_out_csrOp(EX_io_out_csrOp),
    .io_out_takenPre(EX_io_out_takenPre),
    .io_out_takenPrePC(EX_io_out_takenPrePC),
    .io_exeRdData(EX_io_exeRdData),
    .io_bubbleEx(EX_io_bubbleEx),
    .io_takenValid(EX_io_takenValid),
    .io_takenValidJalr(EX_io_takenValidJalr),
    .io_takenMiss(EX_io_takenMiss),
    .io_exTakenPre(EX_io_exTakenPre),
    .io_takenPC(EX_io_takenPC),
    .io_exeX1En(EX_io_exeX1En),
    .io_exeAluRes(EX_io_exeAluRes),
    .io_exc(EX_io_exc),
    .io_csrOp(EX_io_csrOp),
    .io_mepc(EX_io_mepc),
    .io_mtvec(EX_io_mtvec),
    .io_time_int(EX_io_time_int)
  );
  PipelineReg ExRegMem ( // @[Core.scala 21:24]
    .clock(ExRegMem_clock),
    .reset(ExRegMem_reset),
    .io_in_valid(ExRegMem_io_in_valid),
    .io_in_pc(ExRegMem_io_in_pc),
    .io_in_inst(ExRegMem_io_in_inst),
    .io_in_typeL(ExRegMem_io_in_typeL),
    .io_in_aluA(ExRegMem_io_in_aluA),
    .io_in_aluB(ExRegMem_io_in_aluB),
    .io_in_aluOp(ExRegMem_io_in_aluOp),
    .io_in_branch(ExRegMem_io_in_branch),
    .io_in_memtoReg(ExRegMem_io_in_memtoReg),
    .io_in_memWr(ExRegMem_io_in_memWr),
    .io_in_memOp(ExRegMem_io_in_memOp),
    .io_in_memAddr(ExRegMem_io_in_memAddr),
    .io_in_rdEn(ExRegMem_io_in_rdEn),
    .io_in_rdAddr(ExRegMem_io_in_rdAddr),
    .io_in_rs1Data(ExRegMem_io_in_rs1Data),
    .io_in_rs2Data(ExRegMem_io_in_rs2Data),
    .io_in_imm(ExRegMem_io_in_imm),
    .io_in_aluRes(ExRegMem_io_in_aluRes),
    .io_in_memData(ExRegMem_io_in_memData),
    .io_in_csrOp(ExRegMem_io_in_csrOp),
    .io_in_takenPre(ExRegMem_io_in_takenPre),
    .io_in_takenPrePC(ExRegMem_io_in_takenPrePC),
    .io_out_valid(ExRegMem_io_out_valid),
    .io_out_pc(ExRegMem_io_out_pc),
    .io_out_inst(ExRegMem_io_out_inst),
    .io_out_typeL(ExRegMem_io_out_typeL),
    .io_out_aluA(ExRegMem_io_out_aluA),
    .io_out_aluB(ExRegMem_io_out_aluB),
    .io_out_aluOp(ExRegMem_io_out_aluOp),
    .io_out_branch(ExRegMem_io_out_branch),
    .io_out_memtoReg(ExRegMem_io_out_memtoReg),
    .io_out_memWr(ExRegMem_io_out_memWr),
    .io_out_memOp(ExRegMem_io_out_memOp),
    .io_out_memAddr(ExRegMem_io_out_memAddr),
    .io_out_rdEn(ExRegMem_io_out_rdEn),
    .io_out_rdAddr(ExRegMem_io_out_rdAddr),
    .io_out_rs1Data(ExRegMem_io_out_rs1Data),
    .io_out_rs2Data(ExRegMem_io_out_rs2Data),
    .io_out_imm(ExRegMem_io_out_imm),
    .io_out_aluRes(ExRegMem_io_out_aluRes),
    .io_out_memData(ExRegMem_io_out_memData),
    .io_out_csrOp(ExRegMem_io_out_csrOp),
    .io_out_takenPre(ExRegMem_io_out_takenPre),
    .io_out_takenPrePC(ExRegMem_io_out_takenPrePC),
    .io_flush(ExRegMem_io_flush),
    .io_stall(ExRegMem_io_stall)
  );
  DataMem MEM ( // @[Core.scala 22:19]
    .clock(MEM_clock),
    .reset(MEM_reset),
    .io_dmem_data_valid(MEM_io_dmem_data_valid),
    .io_dmem_data_ready(MEM_io_dmem_data_ready),
    .io_dmem_data_req(MEM_io_dmem_data_req),
    .io_dmem_data_addr(MEM_io_dmem_data_addr),
    .io_dmem_data_size(MEM_io_dmem_data_size),
    .io_dmem_data_strb(MEM_io_dmem_data_strb),
    .io_dmem_data_read(MEM_io_dmem_data_read),
    .io_dmem_data_write(MEM_io_dmem_data_write),
    .io_IFDone(MEM_io_IFDone),
    .io_in_valid(MEM_io_in_valid),
    .io_in_pc(MEM_io_in_pc),
    .io_in_inst(MEM_io_in_inst),
    .io_in_typeL(MEM_io_in_typeL),
    .io_in_aluA(MEM_io_in_aluA),
    .io_in_aluB(MEM_io_in_aluB),
    .io_in_aluOp(MEM_io_in_aluOp),
    .io_in_branch(MEM_io_in_branch),
    .io_in_memtoReg(MEM_io_in_memtoReg),
    .io_in_memWr(MEM_io_in_memWr),
    .io_in_memOp(MEM_io_in_memOp),
    .io_in_rdEn(MEM_io_in_rdEn),
    .io_in_rdAddr(MEM_io_in_rdAddr),
    .io_in_rs1Data(MEM_io_in_rs1Data),
    .io_in_rs2Data(MEM_io_in_rs2Data),
    .io_in_imm(MEM_io_in_imm),
    .io_in_aluRes(MEM_io_in_aluRes),
    .io_in_csrOp(MEM_io_in_csrOp),
    .io_in_takenPre(MEM_io_in_takenPre),
    .io_in_takenPrePC(MEM_io_in_takenPrePC),
    .io_out_valid(MEM_io_out_valid),
    .io_out_pc(MEM_io_out_pc),
    .io_out_inst(MEM_io_out_inst),
    .io_out_typeL(MEM_io_out_typeL),
    .io_out_aluA(MEM_io_out_aluA),
    .io_out_aluB(MEM_io_out_aluB),
    .io_out_aluOp(MEM_io_out_aluOp),
    .io_out_branch(MEM_io_out_branch),
    .io_out_memtoReg(MEM_io_out_memtoReg),
    .io_out_memWr(MEM_io_out_memWr),
    .io_out_memOp(MEM_io_out_memOp),
    .io_out_memAddr(MEM_io_out_memAddr),
    .io_out_rdEn(MEM_io_out_rdEn),
    .io_out_rdAddr(MEM_io_out_rdAddr),
    .io_out_rs1Data(MEM_io_out_rs1Data),
    .io_out_rs2Data(MEM_io_out_rs2Data),
    .io_out_imm(MEM_io_out_imm),
    .io_out_aluRes(MEM_io_out_aluRes),
    .io_out_memData(MEM_io_out_memData),
    .io_out_csrOp(MEM_io_out_csrOp),
    .io_out_takenPre(MEM_io_out_takenPre),
    .io_out_takenPrePC(MEM_io_out_takenPrePC),
    .io_memRdData(MEM_io_memRdData),
    .io_memDone(MEM_io_memDone),
    .io_memX1En(MEM_io_memX1En),
    .io_memAluRes(MEM_io_memAluRes),
    .io_cmp_ren(MEM_io_cmp_ren),
    .io_cmp_wen(MEM_io_cmp_wen),
    .io_cmp_addr(MEM_io_cmp_addr),
    .io_cmp_wdata(MEM_io_cmp_wdata),
    .io_cmp_rdata(MEM_io_cmp_rdata)
  );
  PipelineReg MemRegWb ( // @[Core.scala 23:24]
    .clock(MemRegWb_clock),
    .reset(MemRegWb_reset),
    .io_in_valid(MemRegWb_io_in_valid),
    .io_in_pc(MemRegWb_io_in_pc),
    .io_in_inst(MemRegWb_io_in_inst),
    .io_in_typeL(MemRegWb_io_in_typeL),
    .io_in_aluA(MemRegWb_io_in_aluA),
    .io_in_aluB(MemRegWb_io_in_aluB),
    .io_in_aluOp(MemRegWb_io_in_aluOp),
    .io_in_branch(MemRegWb_io_in_branch),
    .io_in_memtoReg(MemRegWb_io_in_memtoReg),
    .io_in_memWr(MemRegWb_io_in_memWr),
    .io_in_memOp(MemRegWb_io_in_memOp),
    .io_in_memAddr(MemRegWb_io_in_memAddr),
    .io_in_rdEn(MemRegWb_io_in_rdEn),
    .io_in_rdAddr(MemRegWb_io_in_rdAddr),
    .io_in_rs1Data(MemRegWb_io_in_rs1Data),
    .io_in_rs2Data(MemRegWb_io_in_rs2Data),
    .io_in_imm(MemRegWb_io_in_imm),
    .io_in_aluRes(MemRegWb_io_in_aluRes),
    .io_in_memData(MemRegWb_io_in_memData),
    .io_in_csrOp(MemRegWb_io_in_csrOp),
    .io_in_takenPre(MemRegWb_io_in_takenPre),
    .io_in_takenPrePC(MemRegWb_io_in_takenPrePC),
    .io_out_valid(MemRegWb_io_out_valid),
    .io_out_pc(MemRegWb_io_out_pc),
    .io_out_inst(MemRegWb_io_out_inst),
    .io_out_typeL(MemRegWb_io_out_typeL),
    .io_out_aluA(MemRegWb_io_out_aluA),
    .io_out_aluB(MemRegWb_io_out_aluB),
    .io_out_aluOp(MemRegWb_io_out_aluOp),
    .io_out_branch(MemRegWb_io_out_branch),
    .io_out_memtoReg(MemRegWb_io_out_memtoReg),
    .io_out_memWr(MemRegWb_io_out_memWr),
    .io_out_memOp(MemRegWb_io_out_memOp),
    .io_out_memAddr(MemRegWb_io_out_memAddr),
    .io_out_rdEn(MemRegWb_io_out_rdEn),
    .io_out_rdAddr(MemRegWb_io_out_rdAddr),
    .io_out_rs1Data(MemRegWb_io_out_rs1Data),
    .io_out_rs2Data(MemRegWb_io_out_rs2Data),
    .io_out_imm(MemRegWb_io_out_imm),
    .io_out_aluRes(MemRegWb_io_out_aluRes),
    .io_out_memData(MemRegWb_io_out_memData),
    .io_out_csrOp(MemRegWb_io_out_csrOp),
    .io_out_takenPre(MemRegWb_io_out_takenPre),
    .io_out_takenPrePC(MemRegWb_io_out_takenPrePC),
    .io_flush(MemRegWb_io_flush),
    .io_stall(MemRegWb_io_stall)
  );
  WriteBack WB ( // @[Core.scala 24:18]
    .clock(WB_clock),
    .reset(WB_reset),
    .io_in_valid(WB_io_in_valid),
    .io_in_pc(WB_io_in_pc),
    .io_in_inst(WB_io_in_inst),
    .io_in_memtoReg(WB_io_in_memtoReg),
    .io_in_memWr(WB_io_in_memWr),
    .io_in_memAddr(WB_io_in_memAddr),
    .io_in_rdEn(WB_io_in_rdEn),
    .io_in_rdAddr(WB_io_in_rdAddr),
    .io_in_rs1Data(WB_io_in_rs1Data),
    .io_in_aluRes(WB_io_in_aluRes),
    .io_in_memData(WB_io_in_memData),
    .io_in_csrOp(WB_io_in_csrOp),
    .io_IFDone(WB_io_IFDone),
    .io_memDone(WB_io_memDone),
    .io_pc_intr(WB_io_pc_intr),
    .io_pc(WB_io_pc),
    .io_inst(WB_io_inst),
    .io_wbRdEn(WB_io_wbRdEn),
    .io_wbRdAddr(WB_io_wbRdAddr),
    .io_wbRdData(WB_io_wbRdData),
    .io_ready_cmt(WB_io_ready_cmt),
    .io_csrOp_WB(WB_io_csrOp_WB),
    .io_mepc(WB_io_mepc),
    .io_mtvec(WB_io_mtvec),
    .io_cmp_ren(WB_io_cmp_ren),
    .io_cmp_wen(WB_io_cmp_wen),
    .io_cmp_addr(WB_io_cmp_addr),
    .io_cmp_wdata(WB_io_cmp_wdata),
    .io_cmp_rdata(WB_io_cmp_rdata),
    .io_exc(WB_io_exc),
    .io_memtoReg(WB_io_memtoReg),
    .io_memWr(WB_io_memWr),
    .io_mem_addr(WB_io_mem_addr),
    .io_time_int(WB_io_time_int)
  );
  preDebug preDebug ( // @[Core.scala 27:24]
    .clock(preDebug_clock),
    .reset(preDebug_reset),
    .io_exeBranch(preDebug_io_exeBranch),
    .io_takenMiss(preDebug_io_takenMiss),
    .io_rs1Addr(preDebug_io_rs1Addr),
    .io_coreEnd(preDebug_io_coreEnd),
    .io_IFDone(preDebug_io_IFDone),
    .io_memDone(preDebug_io_memDone)
  );
  DifftestInstrCommit dt_ic ( // @[Core.scala 166:21]
    .clock(dt_ic_clock),
    .coreid(dt_ic_coreid),
    .index(dt_ic_index),
    .valid(dt_ic_valid),
    .pc(dt_ic_pc),
    .instr(dt_ic_instr),
    .skip(dt_ic_skip),
    .isRVC(dt_ic_isRVC),
    .scFailed(dt_ic_scFailed),
    .wen(dt_ic_wen),
    .wdata(dt_ic_wdata),
    .wdest(dt_ic_wdest)
  );
  DifftestArchEvent dt_ae ( // @[Core.scala 180:21]
    .clock(dt_ae_clock),
    .coreid(dt_ae_coreid),
    .intrNO(dt_ae_intrNO),
    .cause(dt_ae_cause),
    .exceptionPC(dt_ae_exceptionPC),
    .exceptionInst(dt_ae_exceptionInst)
  );
  DifftestTrapEvent dt_te ( // @[Core.scala 193:21]
    .clock(dt_te_clock),
    .coreid(dt_te_coreid),
    .valid(dt_te_valid),
    .code(dt_te_code),
    .pc(dt_te_pc),
    .cycleCnt(dt_te_cycleCnt),
    .instrCnt(dt_te_instrCnt)
  );
  assign io_imem_inst_valid = IF_io_imem_inst_valid; // @[Core.scala 66:22]
  assign io_imem_inst_addr = IF_io_imem_inst_addr; // @[Core.scala 68:21]
  assign io_dmem_data_valid = MEM_io_dmem_data_valid; // @[Core.scala 135:15]
  assign io_dmem_data_req = MEM_io_dmem_data_req; // @[Core.scala 135:15]
  assign io_dmem_data_addr = MEM_io_dmem_data_addr; // @[Core.scala 135:15]
  assign io_dmem_data_size = MEM_io_dmem_data_size; // @[Core.scala 135:15]
  assign io_dmem_data_strb = MEM_io_dmem_data_strb; // @[Core.scala 135:15]
  assign io_dmem_data_write = MEM_io_dmem_data_write; // @[Core.scala 135:15]
  assign IF_clock = clock;
  assign IF_reset = reset;
  assign IF_io_imem_inst_ready = io_imem_inst_ready; // @[Core.scala 72:25]
  assign IF_io_imem_inst_read = io_imem_inst_read; // @[Core.scala 71:24]
  assign IF_io_takenValid = EX_io_takenValid; // @[Core.scala 74:20]
  assign IF_io_takenValidJalr = EX_io_takenValidJalr; // @[Core.scala 75:24]
  assign IF_io_takenMiss = EX_io_takenMiss; // @[Core.scala 76:19]
  assign IF_io_exTakenPre = EX_io_exTakenPre; // @[Core.scala 77:20]
  assign IF_io_takenPC = EX_io_takenPC; // @[Core.scala 78:17]
  assign IF_io_nextPC = EX_io_out_nextPC; // @[Core.scala 79:16]
  assign IF_io_stall = EXLHitID | _stallIfIdEn_T_1 | EXSHitIDEn; // @[Core.scala 91:46]
  assign IF_io_exc = WB_io_exc; // @[Core.scala 92:13]
  assign IF_io_intr = WB_io_time_int; // @[Core.scala 93:14]
  assign IF_io_preRs1Data = ID_io_preRs1Data; // @[Core.scala 81:20]
  assign IF_io_preRs1x1Data = ID_io_preRs1x1Data; // @[Core.scala 82:22]
  assign IF_io_exeX1En = EX_io_exeX1En; // @[Core.scala 83:17]
  assign IF_io_exeAluRes = EX_io_exeAluRes; // @[Core.scala 84:19]
  assign IF_io_memX1En = MEM_io_memX1En; // @[Core.scala 85:17]
  assign IF_io_memAluRes = MEM_io_memAluRes; // @[Core.scala 86:19]
  assign IF_io_wbRdEn = WB_io_wbRdEn; // @[Core.scala 87:16]
  assign IF_io_wbRdAddr = WB_io_wbRdAddr; // @[Core.scala 88:18]
  assign IF_io_wbRdData = WB_io_wbRdData; // @[Core.scala 89:18]
  assign IfRegId_clock = clock;
  assign IfRegId_reset = reset;
  assign IfRegId_io_in_valid = IF_io_out_valid; // @[Core.scala 95:17]
  assign IfRegId_io_in_pc = IF_io_out_pc; // @[Core.scala 95:17]
  assign IfRegId_io_in_inst = IF_io_out_inst; // @[Core.scala 95:17]
  assign IfRegId_io_in_typeL = 1'h0; // @[Core.scala 95:17]
  assign IfRegId_io_in_aluA = 1'h0; // @[Core.scala 95:17]
  assign IfRegId_io_in_aluB = 2'h0; // @[Core.scala 95:17]
  assign IfRegId_io_in_aluOp = 4'h0; // @[Core.scala 95:17]
  assign IfRegId_io_in_branch = 3'h0; // @[Core.scala 95:17]
  assign IfRegId_io_in_memtoReg = 2'h0; // @[Core.scala 95:17]
  assign IfRegId_io_in_memWr = 1'h0; // @[Core.scala 95:17]
  assign IfRegId_io_in_memOp = 3'h0; // @[Core.scala 95:17]
  assign IfRegId_io_in_memAddr = 32'h0; // @[Core.scala 95:17]
  assign IfRegId_io_in_rdEn = 1'h0; // @[Core.scala 95:17]
  assign IfRegId_io_in_rdAddr = 5'h0; // @[Core.scala 95:17]
  assign IfRegId_io_in_rs1Data = 64'h0; // @[Core.scala 95:17]
  assign IfRegId_io_in_rs2Data = 64'h0; // @[Core.scala 95:17]
  assign IfRegId_io_in_imm = 64'h0; // @[Core.scala 95:17]
  assign IfRegId_io_in_aluRes = 64'h0; // @[Core.scala 95:17]
  assign IfRegId_io_in_memData = 64'h0; // @[Core.scala 95:17]
  assign IfRegId_io_in_csrOp = 4'h0; // @[Core.scala 95:17]
  assign IfRegId_io_in_takenPre = IF_io_out_takenPre; // @[Core.scala 95:17]
  assign IfRegId_io_in_takenPrePC = IF_io_out_takenPrePC; // @[Core.scala 95:17]
  assign IfRegId_io_flush = ecallEn | WB_io_time_int | EX_io_takenMiss; // @[Core.scala 51:38]
  assign IfRegId_io_stall = ~IF_io_IFDone | ~MEM_io_memDone | (EXLHitID | EXSHitIDEn) & ~WB_io_time_int; // @[Core.scala 59:55]
  assign ID_clock = clock;
  assign ID_reset = reset;
  assign ID_io_rdEn = WB_io_wbRdEn; // @[Core.scala 100:14]
  assign ID_io_rdAddr = WB_io_wbRdAddr; // @[Core.scala 101:16]
  assign ID_io_rdData = WB_io_wbRdData; // @[Core.scala 102:16]
  assign ID_io_preRs1En = IF_io_preRs1En; // @[Core.scala 104:18]
  assign ID_io_preRs1Addr = IF_io_preRs1Addr; // @[Core.scala 105:20]
  assign ID_io_in_valid = IfRegId_io_out_valid; // @[Core.scala 99:12]
  assign ID_io_in_pc = IfRegId_io_out_pc; // @[Core.scala 99:12]
  assign ID_io_in_inst = IfRegId_io_out_inst; // @[Core.scala 99:12]
  assign ID_io_in_takenPre = IfRegId_io_out_takenPre; // @[Core.scala 99:12]
  assign ID_io_in_takenPrePC = IfRegId_io_out_takenPrePC; // @[Core.scala 99:12]
  assign ID_io_exeRdEn = EX_io_out_rdEn; // @[Core.scala 107:17]
  assign ID_io_exeRdAddr = EX_io_out_rdAddr; // @[Core.scala 108:19]
  assign ID_io_exeRdData = EX_io_exeRdData; // @[Core.scala 109:19]
  assign ID_io_memRdEn = MEM_io_out_rdEn; // @[Core.scala 111:17]
  assign ID_io_memRdAddr = MEM_io_out_rdAddr; // @[Core.scala 112:19]
  assign ID_io_memRdData = MEM_io_memRdData; // @[Core.scala 113:19]
  assign ID_io_wbRdEn = WB_io_wbRdEn; // @[Core.scala 115:16]
  assign ID_io_wbRdAddr = WB_io_wbRdAddr; // @[Core.scala 116:18]
  assign ID_io_wbRdData = WB_io_wbRdData; // @[Core.scala 117:18]
  assign IdRegEx_clock = clock;
  assign IdRegEx_reset = reset;
  assign IdRegEx_io_in_valid = ID_io_out_valid; // @[Core.scala 119:17]
  assign IdRegEx_io_in_pc = ID_io_out_pc; // @[Core.scala 119:17]
  assign IdRegEx_io_in_inst = ID_io_out_inst; // @[Core.scala 119:17]
  assign IdRegEx_io_in_typeL = ID_io_out_typeL; // @[Core.scala 119:17]
  assign IdRegEx_io_in_aluA = ID_io_out_aluA; // @[Core.scala 119:17]
  assign IdRegEx_io_in_aluB = ID_io_out_aluB; // @[Core.scala 119:17]
  assign IdRegEx_io_in_aluOp = ID_io_out_aluOp; // @[Core.scala 119:17]
  assign IdRegEx_io_in_branch = ID_io_out_branch; // @[Core.scala 119:17]
  assign IdRegEx_io_in_memtoReg = ID_io_out_memtoReg; // @[Core.scala 119:17]
  assign IdRegEx_io_in_memWr = ID_io_out_memWr; // @[Core.scala 119:17]
  assign IdRegEx_io_in_memOp = ID_io_out_memOp; // @[Core.scala 119:17]
  assign IdRegEx_io_in_memAddr = 32'h0; // @[Core.scala 119:17]
  assign IdRegEx_io_in_rdEn = ID_io_out_rdEn; // @[Core.scala 119:17]
  assign IdRegEx_io_in_rdAddr = ID_io_out_rdAddr; // @[Core.scala 119:17]
  assign IdRegEx_io_in_rs1Data = ID_io_out_rs1Data; // @[Core.scala 119:17]
  assign IdRegEx_io_in_rs2Data = ID_io_out_rs2Data; // @[Core.scala 119:17]
  assign IdRegEx_io_in_imm = ID_io_out_imm; // @[Core.scala 119:17]
  assign IdRegEx_io_in_aluRes = 64'h0; // @[Core.scala 119:17]
  assign IdRegEx_io_in_memData = 64'h0; // @[Core.scala 119:17]
  assign IdRegEx_io_in_csrOp = ID_io_out_csrOp; // @[Core.scala 119:17]
  assign IdRegEx_io_in_takenPre = ID_io_out_takenPre; // @[Core.scala 119:17]
  assign IdRegEx_io_in_takenPrePC = ID_io_out_takenPrePC; // @[Core.scala 119:17]
  assign IdRegEx_io_flush = ecallEn | IF_io_IFDone & (EX_io_takenMiss | EXLHitID | EXSHitIDEn); // @[Core.scala 52:25]
  assign IdRegEx_io_stall = _stallIfIdEn_T | _stallIfIdEn_T_1; // @[Core.scala 60:36]
  assign EX_io_in_valid = IdRegEx_io_out_valid; // @[Core.scala 123:12]
  assign EX_io_in_pc = IdRegEx_io_out_pc; // @[Core.scala 123:12]
  assign EX_io_in_inst = IdRegEx_io_out_inst; // @[Core.scala 123:12]
  assign EX_io_in_typeL = IdRegEx_io_out_typeL; // @[Core.scala 123:12]
  assign EX_io_in_aluA = IdRegEx_io_out_aluA; // @[Core.scala 123:12]
  assign EX_io_in_aluB = IdRegEx_io_out_aluB; // @[Core.scala 123:12]
  assign EX_io_in_aluOp = IdRegEx_io_out_aluOp; // @[Core.scala 123:12]
  assign EX_io_in_branch = IdRegEx_io_out_branch; // @[Core.scala 123:12]
  assign EX_io_in_memtoReg = IdRegEx_io_out_memtoReg; // @[Core.scala 123:12]
  assign EX_io_in_memWr = IdRegEx_io_out_memWr; // @[Core.scala 123:12]
  assign EX_io_in_memOp = IdRegEx_io_out_memOp; // @[Core.scala 123:12]
  assign EX_io_in_rdEn = IdRegEx_io_out_rdEn; // @[Core.scala 123:12]
  assign EX_io_in_rdAddr = IdRegEx_io_out_rdAddr; // @[Core.scala 123:12]
  assign EX_io_in_rs1Data = IdRegEx_io_out_rs1Data; // @[Core.scala 123:12]
  assign EX_io_in_rs2Data = IdRegEx_io_out_rs2Data; // @[Core.scala 123:12]
  assign EX_io_in_imm = IdRegEx_io_out_imm; // @[Core.scala 123:12]
  assign EX_io_in_csrOp = IdRegEx_io_out_csrOp; // @[Core.scala 123:12]
  assign EX_io_in_takenPre = IdRegEx_io_out_takenPre; // @[Core.scala 123:12]
  assign EX_io_in_takenPrePC = IdRegEx_io_out_takenPrePC; // @[Core.scala 123:12]
  assign EX_io_exc = WB_io_exc; // @[Core.scala 124:13]
  assign EX_io_csrOp = WB_io_csrOp_WB; // @[Core.scala 125:15]
  assign EX_io_mepc = WB_io_mepc; // @[Core.scala 126:14]
  assign EX_io_mtvec = WB_io_mtvec; // @[Core.scala 127:15]
  assign EX_io_time_int = WB_io_time_int; // @[Core.scala 128:18]
  assign ExRegMem_clock = clock;
  assign ExRegMem_reset = reset;
  assign ExRegMem_io_in_valid = EX_io_out_valid; // @[Core.scala 130:18]
  assign ExRegMem_io_in_pc = EX_io_out_pc; // @[Core.scala 130:18]
  assign ExRegMem_io_in_inst = EX_io_out_inst; // @[Core.scala 130:18]
  assign ExRegMem_io_in_typeL = EX_io_out_typeL; // @[Core.scala 130:18]
  assign ExRegMem_io_in_aluA = EX_io_out_aluA; // @[Core.scala 130:18]
  assign ExRegMem_io_in_aluB = EX_io_out_aluB; // @[Core.scala 130:18]
  assign ExRegMem_io_in_aluOp = EX_io_out_aluOp; // @[Core.scala 130:18]
  assign ExRegMem_io_in_branch = EX_io_out_branch; // @[Core.scala 130:18]
  assign ExRegMem_io_in_memtoReg = EX_io_out_memtoReg; // @[Core.scala 130:18]
  assign ExRegMem_io_in_memWr = EX_io_out_memWr; // @[Core.scala 130:18]
  assign ExRegMem_io_in_memOp = EX_io_out_memOp; // @[Core.scala 130:18]
  assign ExRegMem_io_in_memAddr = 32'h0; // @[Core.scala 130:18]
  assign ExRegMem_io_in_rdEn = EX_io_out_rdEn; // @[Core.scala 130:18]
  assign ExRegMem_io_in_rdAddr = EX_io_out_rdAddr; // @[Core.scala 130:18]
  assign ExRegMem_io_in_rs1Data = EX_io_out_rs1Data; // @[Core.scala 130:18]
  assign ExRegMem_io_in_rs2Data = EX_io_out_rs2Data; // @[Core.scala 130:18]
  assign ExRegMem_io_in_imm = EX_io_out_imm; // @[Core.scala 130:18]
  assign ExRegMem_io_in_aluRes = EX_io_out_aluRes; // @[Core.scala 130:18]
  assign ExRegMem_io_in_memData = 64'h0; // @[Core.scala 130:18]
  assign ExRegMem_io_in_csrOp = EX_io_out_csrOp; // @[Core.scala 130:18]
  assign ExRegMem_io_in_takenPre = EX_io_out_takenPre; // @[Core.scala 130:18]
  assign ExRegMem_io_in_takenPrePC = EX_io_out_takenPrePC; // @[Core.scala 130:18]
  assign ExRegMem_io_flush = WB_io_csrOp_WB[3] | WB_io_time_int; // @[Core.scala 50:43]
  assign ExRegMem_io_stall = _stallIfIdEn_T | _stallIfIdEn_T_1; // @[Core.scala 61:36]
  assign MEM_clock = clock;
  assign MEM_reset = reset;
  assign MEM_io_dmem_data_ready = io_dmem_data_ready; // @[Core.scala 135:15]
  assign MEM_io_dmem_data_read = io_dmem_data_read; // @[Core.scala 135:15]
  assign MEM_io_IFDone = IF_io_IFDone; // @[Core.scala 136:17]
  assign MEM_io_in_valid = ExRegMem_io_out_valid; // @[Core.scala 134:13]
  assign MEM_io_in_pc = ExRegMem_io_out_pc; // @[Core.scala 134:13]
  assign MEM_io_in_inst = ExRegMem_io_out_inst; // @[Core.scala 134:13]
  assign MEM_io_in_typeL = ExRegMem_io_out_typeL; // @[Core.scala 134:13]
  assign MEM_io_in_aluA = ExRegMem_io_out_aluA; // @[Core.scala 134:13]
  assign MEM_io_in_aluB = ExRegMem_io_out_aluB; // @[Core.scala 134:13]
  assign MEM_io_in_aluOp = ExRegMem_io_out_aluOp; // @[Core.scala 134:13]
  assign MEM_io_in_branch = ExRegMem_io_out_branch; // @[Core.scala 134:13]
  assign MEM_io_in_memtoReg = ExRegMem_io_out_memtoReg; // @[Core.scala 134:13]
  assign MEM_io_in_memWr = ExRegMem_io_out_memWr; // @[Core.scala 134:13]
  assign MEM_io_in_memOp = ExRegMem_io_out_memOp; // @[Core.scala 134:13]
  assign MEM_io_in_rdEn = ExRegMem_io_out_rdEn; // @[Core.scala 134:13]
  assign MEM_io_in_rdAddr = ExRegMem_io_out_rdAddr; // @[Core.scala 134:13]
  assign MEM_io_in_rs1Data = ExRegMem_io_out_rs1Data; // @[Core.scala 134:13]
  assign MEM_io_in_rs2Data = ExRegMem_io_out_rs2Data; // @[Core.scala 134:13]
  assign MEM_io_in_imm = ExRegMem_io_out_imm; // @[Core.scala 134:13]
  assign MEM_io_in_aluRes = ExRegMem_io_out_aluRes; // @[Core.scala 134:13]
  assign MEM_io_in_csrOp = ExRegMem_io_out_csrOp; // @[Core.scala 134:13]
  assign MEM_io_in_takenPre = ExRegMem_io_out_takenPre; // @[Core.scala 134:13]
  assign MEM_io_in_takenPrePC = ExRegMem_io_out_takenPrePC; // @[Core.scala 134:13]
  assign MEM_io_cmp_rdata = WB_io_cmp_rdata; // @[Core.scala 137:20]
  assign MemRegWb_clock = clock;
  assign MemRegWb_reset = reset;
  assign MemRegWb_io_in_valid = MEM_io_out_valid; // @[Core.scala 139:18]
  assign MemRegWb_io_in_pc = MEM_io_out_pc; // @[Core.scala 139:18]
  assign MemRegWb_io_in_inst = MEM_io_out_inst; // @[Core.scala 139:18]
  assign MemRegWb_io_in_typeL = MEM_io_out_typeL; // @[Core.scala 139:18]
  assign MemRegWb_io_in_aluA = MEM_io_out_aluA; // @[Core.scala 139:18]
  assign MemRegWb_io_in_aluB = MEM_io_out_aluB; // @[Core.scala 139:18]
  assign MemRegWb_io_in_aluOp = MEM_io_out_aluOp; // @[Core.scala 139:18]
  assign MemRegWb_io_in_branch = MEM_io_out_branch; // @[Core.scala 139:18]
  assign MemRegWb_io_in_memtoReg = MEM_io_out_memtoReg; // @[Core.scala 139:18]
  assign MemRegWb_io_in_memWr = MEM_io_out_memWr; // @[Core.scala 139:18]
  assign MemRegWb_io_in_memOp = MEM_io_out_memOp; // @[Core.scala 139:18]
  assign MemRegWb_io_in_memAddr = MEM_io_out_memAddr; // @[Core.scala 139:18]
  assign MemRegWb_io_in_rdEn = MEM_io_out_rdEn; // @[Core.scala 139:18]
  assign MemRegWb_io_in_rdAddr = MEM_io_out_rdAddr; // @[Core.scala 139:18]
  assign MemRegWb_io_in_rs1Data = MEM_io_out_rs1Data; // @[Core.scala 139:18]
  assign MemRegWb_io_in_rs2Data = MEM_io_out_rs2Data; // @[Core.scala 139:18]
  assign MemRegWb_io_in_imm = MEM_io_out_imm; // @[Core.scala 139:18]
  assign MemRegWb_io_in_aluRes = MEM_io_out_aluRes; // @[Core.scala 139:18]
  assign MemRegWb_io_in_memData = MEM_io_out_memData; // @[Core.scala 139:18]
  assign MemRegWb_io_in_csrOp = MEM_io_out_csrOp; // @[Core.scala 139:18]
  assign MemRegWb_io_in_takenPre = MEM_io_out_takenPre; // @[Core.scala 139:18]
  assign MemRegWb_io_in_takenPrePC = MEM_io_out_takenPrePC; // @[Core.scala 139:18]
  assign MemRegWb_io_flush = WB_io_csrOp_WB[3] | WB_io_time_int; // @[Core.scala 50:43]
  assign MemRegWb_io_stall = _stallIfIdEn_T | _stallIfIdEn_T_1; // @[Core.scala 62:36]
  assign WB_clock = clock;
  assign WB_reset = reset;
  assign WB_io_in_valid = MemRegWb_io_out_valid; // @[Core.scala 143:12]
  assign WB_io_in_pc = MemRegWb_io_out_pc; // @[Core.scala 143:12]
  assign WB_io_in_inst = MemRegWb_io_out_inst; // @[Core.scala 143:12]
  assign WB_io_in_memtoReg = MemRegWb_io_out_memtoReg; // @[Core.scala 143:12]
  assign WB_io_in_memWr = MemRegWb_io_out_memWr; // @[Core.scala 143:12]
  assign WB_io_in_memAddr = MemRegWb_io_out_memAddr; // @[Core.scala 143:12]
  assign WB_io_in_rdEn = MemRegWb_io_out_rdEn; // @[Core.scala 143:12]
  assign WB_io_in_rdAddr = MemRegWb_io_out_rdAddr; // @[Core.scala 143:12]
  assign WB_io_in_rs1Data = MemRegWb_io_out_rs1Data; // @[Core.scala 143:12]
  assign WB_io_in_aluRes = MemRegWb_io_out_aluRes; // @[Core.scala 143:12]
  assign WB_io_in_memData = MemRegWb_io_out_memData; // @[Core.scala 143:12]
  assign WB_io_in_csrOp = MemRegWb_io_out_csrOp; // @[Core.scala 143:12]
  assign WB_io_IFDone = IF_io_IFDone; // @[Core.scala 144:16]
  assign WB_io_memDone = MEM_io_memDone; // @[Core.scala 145:17]
  assign WB_io_pc_intr = WB_io_time_int ? _exceptionPC_T_7 : 32'h0; // @[Core.scala 37:24]
  assign WB_io_cmp_ren = MEM_io_cmp_ren; // @[Core.scala 147:17]
  assign WB_io_cmp_wen = MEM_io_cmp_wen; // @[Core.scala 148:17]
  assign WB_io_cmp_addr = MEM_io_cmp_addr; // @[Core.scala 149:18]
  assign WB_io_cmp_wdata = MEM_io_cmp_wdata; // @[Core.scala 150:19]
  assign preDebug_clock = clock;
  assign preDebug_reset = reset;
  assign preDebug_io_exeBranch = EX_io_out_branch; // @[Core.scala 28:25]
  assign preDebug_io_takenMiss = EX_io_takenMiss; // @[Core.scala 29:25]
  assign preDebug_io_rs1Addr = EX_io_out_inst[19:15]; // @[Core.scala 30:40]
  assign preDebug_io_coreEnd = WB_io_inst == 32'h6b; // @[Core.scala 31:37]
  assign preDebug_io_IFDone = IF_io_IFDone; // @[Core.scala 32:22]
  assign preDebug_io_memDone = MEM_io_memDone; // @[Core.scala 33:23]
  assign dt_ic_clock = clock; // @[Core.scala 167:21]
  assign dt_ic_coreid = 8'h0; // @[Core.scala 168:21]
  assign dt_ic_index = 8'h0; // @[Core.scala 169:21]
  assign dt_ic_valid = dt_ic_io_valid_REG; // @[Core.scala 170:21]
  assign dt_ic_pc = {{32'd0}, dt_ic_io_pc_REG}; // @[Core.scala 171:21]
  assign dt_ic_instr = dt_ic_io_instr_REG; // @[Core.scala 172:21]
  assign dt_ic_skip = dt_ic_io_skip_REG; // @[Core.scala 173:21]
  assign dt_ic_isRVC = 1'h0; // @[Core.scala 174:21]
  assign dt_ic_scFailed = 1'h0; // @[Core.scala 175:21]
  assign dt_ic_wen = dt_ic_io_wen_REG; // @[Core.scala 176:21]
  assign dt_ic_wdata = dt_ic_io_wdata_REG; // @[Core.scala 177:21]
  assign dt_ic_wdest = {{3'd0}, dt_ic_io_wdest_REG}; // @[Core.scala 178:21]
  assign dt_ae_clock = clock; // @[Core.scala 181:25]
  assign dt_ae_coreid = 8'h0; // @[Core.scala 182:25]
  assign dt_ae_intrNO = {{29'd0}, dt_ae_io_intrNO_REG}; // @[Core.scala 183:25]
  assign dt_ae_cause = 32'h0; // @[Core.scala 184:25]
  assign dt_ae_exceptionPC = {{32'd0}, dt_ae_io_exceptionPC_REG}; // @[Core.scala 185:25]
  assign dt_ae_exceptionInst = 32'h0;
  assign dt_te_clock = clock; // @[Core.scala 194:21]
  assign dt_te_coreid = 8'h0; // @[Core.scala 195:21]
  assign dt_te_valid = WB_io_inst == 32'h6b; // @[Core.scala 196:36]
  assign dt_te_code = rf_a0_0[2:0]; // @[Core.scala 197:29]
  assign dt_te_pc = {{32'd0}, WB_io_pc}; // @[Core.scala 198:21]
  assign dt_te_cycleCnt = cycle_cnt; // @[Core.scala 199:21]
  assign dt_te_instrCnt = instr_cnt; // @[Core.scala 200:21]
  always @(posedge clock) begin
    dt_ic_io_valid_REG <= WB_io_ready_cmt & IF_io_IFDone & MEM_io_memDone; // @[Core.scala 153:47]
    dt_ic_io_pc_REG <= WB_io_pc; // @[Core.scala 171:31]
    dt_ic_io_instr_REG <= WB_io_inst; // @[Core.scala 172:31]
    dt_ic_io_skip_REG <= _T_1 | WB_io_inst[31:20] == 12'hb00 & WB_io_csrOp_WB != 4'h0 | req_clint; // @[Core.scala 164:102]
    dt_ic_io_wen_REG <= WB_io_wbRdEn; // @[Core.scala 176:31]
    dt_ic_io_wdata_REG <= WB_io_wbRdData; // @[Core.scala 177:31]
    dt_ic_io_wdest_REG <= WB_io_wbRdAddr; // @[Core.scala 178:31]
    if (WB_io_time_int) begin // @[Core.scala 36:20]
      dt_ae_io_intrNO_REG <= 3'h7;
    end else begin
      dt_ae_io_intrNO_REG <= 3'h0;
    end
    if (WB_io_time_int) begin // @[Core.scala 37:24]
      if (WB_io_pc != 32'h0) begin // @[Core.scala 37:34]
        dt_ae_io_exceptionPC_REG <= WB_io_pc;
      end else if (MEM_io_out_pc != 32'h0) begin // @[Core.scala 38:36]
        dt_ae_io_exceptionPC_REG <= MEM_io_out_pc;
      end else if (EX_io_out_pc != 32'h0) begin // @[Core.scala 39:38]
        dt_ae_io_exceptionPC_REG <= EX_io_out_pc;
      end else begin
        dt_ae_io_exceptionPC_REG <= _exceptionPC_T_4;
      end
    end else begin
      dt_ae_io_exceptionPC_REG <= 32'h0;
    end
    if (reset) begin // @[Core.scala 187:26]
      cycle_cnt <= 64'h0; // @[Core.scala 187:26]
    end else begin
      cycle_cnt <= _cycle_cnt_T_1; // @[Core.scala 190:13]
    end
    if (reset) begin // @[Core.scala 188:26]
      instr_cnt <= 64'h0; // @[Core.scala 188:26]
    end else begin
      instr_cnt <= _instr_cnt_T_1; // @[Core.scala 191:13]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~reset) begin
          $fwrite(32'h80000002,"%c",rf_a0_0); // @[Core.scala 159:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  dt_ic_io_valid_REG = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  dt_ic_io_pc_REG = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  dt_ic_io_instr_REG = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  dt_ic_io_skip_REG = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  dt_ic_io_wen_REG = _RAND_4[0:0];
  _RAND_5 = {2{`RANDOM}};
  dt_ic_io_wdata_REG = _RAND_5[63:0];
  _RAND_6 = {1{`RANDOM}};
  dt_ic_io_wdest_REG = _RAND_6[4:0];
  _RAND_7 = {1{`RANDOM}};
  dt_ae_io_intrNO_REG = _RAND_7[2:0];
  _RAND_8 = {1{`RANDOM}};
  dt_ae_io_exceptionPC_REG = _RAND_8[31:0];
  _RAND_9 = {2{`RANDOM}};
  cycle_cnt = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  instr_cnt = _RAND_10[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ICache(
  input          clock,
  input          reset,
  input          io_imem_inst_valid,
  output         io_imem_inst_ready,
  input  [31:0]  io_imem_inst_addr,
  output [31:0]  io_imem_inst_read,
  output         io_out_inst_valid,
  input          io_out_inst_ready,
  output [31:0]  io_out_inst_addr,
  input  [127:0] io_out_inst_read
);
`ifdef RANDOMIZE_REG_INIT
  reg [127:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_645;
  reg [31:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_649;
  reg [31:0] _RAND_650;
  reg [31:0] _RAND_651;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
  reg [31:0] _RAND_654;
  reg [31:0] _RAND_655;
  reg [31:0] _RAND_656;
  reg [31:0] _RAND_657;
  reg [31:0] _RAND_658;
  reg [31:0] _RAND_659;
  reg [31:0] _RAND_660;
  reg [31:0] _RAND_661;
  reg [31:0] _RAND_662;
  reg [31:0] _RAND_663;
  reg [31:0] _RAND_664;
  reg [31:0] _RAND_665;
  reg [31:0] _RAND_666;
  reg [31:0] _RAND_667;
  reg [31:0] _RAND_668;
  reg [31:0] _RAND_669;
  reg [31:0] _RAND_670;
  reg [31:0] _RAND_671;
  reg [31:0] _RAND_672;
  reg [31:0] _RAND_673;
  reg [31:0] _RAND_674;
  reg [31:0] _RAND_675;
  reg [31:0] _RAND_676;
  reg [31:0] _RAND_677;
  reg [31:0] _RAND_678;
  reg [31:0] _RAND_679;
  reg [31:0] _RAND_680;
  reg [31:0] _RAND_681;
  reg [31:0] _RAND_682;
  reg [31:0] _RAND_683;
  reg [31:0] _RAND_684;
  reg [31:0] _RAND_685;
  reg [31:0] _RAND_686;
  reg [31:0] _RAND_687;
  reg [31:0] _RAND_688;
  reg [31:0] _RAND_689;
  reg [31:0] _RAND_690;
  reg [31:0] _RAND_691;
  reg [31:0] _RAND_692;
  reg [31:0] _RAND_693;
  reg [31:0] _RAND_694;
  reg [31:0] _RAND_695;
  reg [31:0] _RAND_696;
  reg [31:0] _RAND_697;
  reg [31:0] _RAND_698;
  reg [31:0] _RAND_699;
  reg [31:0] _RAND_700;
  reg [31:0] _RAND_701;
  reg [31:0] _RAND_702;
  reg [31:0] _RAND_703;
  reg [31:0] _RAND_704;
  reg [31:0] _RAND_705;
  reg [31:0] _RAND_706;
  reg [31:0] _RAND_707;
  reg [31:0] _RAND_708;
  reg [31:0] _RAND_709;
  reg [31:0] _RAND_710;
  reg [31:0] _RAND_711;
  reg [31:0] _RAND_712;
  reg [31:0] _RAND_713;
  reg [31:0] _RAND_714;
  reg [31:0] _RAND_715;
  reg [31:0] _RAND_716;
  reg [31:0] _RAND_717;
  reg [31:0] _RAND_718;
  reg [31:0] _RAND_719;
  reg [31:0] _RAND_720;
  reg [31:0] _RAND_721;
  reg [31:0] _RAND_722;
  reg [31:0] _RAND_723;
  reg [31:0] _RAND_724;
  reg [31:0] _RAND_725;
  reg [31:0] _RAND_726;
  reg [31:0] _RAND_727;
  reg [31:0] _RAND_728;
  reg [31:0] _RAND_729;
  reg [31:0] _RAND_730;
  reg [31:0] _RAND_731;
  reg [31:0] _RAND_732;
  reg [31:0] _RAND_733;
  reg [31:0] _RAND_734;
  reg [31:0] _RAND_735;
  reg [31:0] _RAND_736;
  reg [31:0] _RAND_737;
  reg [31:0] _RAND_738;
  reg [31:0] _RAND_739;
  reg [31:0] _RAND_740;
  reg [31:0] _RAND_741;
  reg [31:0] _RAND_742;
  reg [31:0] _RAND_743;
  reg [31:0] _RAND_744;
  reg [31:0] _RAND_745;
  reg [31:0] _RAND_746;
  reg [31:0] _RAND_747;
  reg [31:0] _RAND_748;
  reg [31:0] _RAND_749;
  reg [31:0] _RAND_750;
  reg [31:0] _RAND_751;
  reg [31:0] _RAND_752;
  reg [31:0] _RAND_753;
  reg [31:0] _RAND_754;
  reg [31:0] _RAND_755;
  reg [31:0] _RAND_756;
  reg [31:0] _RAND_757;
  reg [31:0] _RAND_758;
  reg [31:0] _RAND_759;
  reg [31:0] _RAND_760;
  reg [31:0] _RAND_761;
  reg [31:0] _RAND_762;
  reg [31:0] _RAND_763;
  reg [31:0] _RAND_764;
  reg [31:0] _RAND_765;
  reg [31:0] _RAND_766;
  reg [31:0] _RAND_767;
  reg [31:0] _RAND_768;
  reg [31:0] _RAND_769;
`endif // RANDOMIZE_REG_INIT
  wire [127:0] req_Q; // @[ICache.scala 54:19]
  wire  req_CLK; // @[ICache.scala 54:19]
  wire  req_CEN; // @[ICache.scala 54:19]
  wire  req_WEN; // @[ICache.scala 54:19]
  wire [7:0] req_A; // @[ICache.scala 54:19]
  wire [127:0] req_D; // @[ICache.scala 54:19]
  reg [127:0] cacheWData; // @[ICache.scala 22:27]
  reg  way0V_0; // @[ICache.scala 27:22]
  reg  way0V_1; // @[ICache.scala 27:22]
  reg  way0V_2; // @[ICache.scala 27:22]
  reg  way0V_3; // @[ICache.scala 27:22]
  reg  way0V_4; // @[ICache.scala 27:22]
  reg  way0V_5; // @[ICache.scala 27:22]
  reg  way0V_6; // @[ICache.scala 27:22]
  reg  way0V_7; // @[ICache.scala 27:22]
  reg  way0V_8; // @[ICache.scala 27:22]
  reg  way0V_9; // @[ICache.scala 27:22]
  reg  way0V_10; // @[ICache.scala 27:22]
  reg  way0V_11; // @[ICache.scala 27:22]
  reg  way0V_12; // @[ICache.scala 27:22]
  reg  way0V_13; // @[ICache.scala 27:22]
  reg  way0V_14; // @[ICache.scala 27:22]
  reg  way0V_15; // @[ICache.scala 27:22]
  reg  way0V_16; // @[ICache.scala 27:22]
  reg  way0V_17; // @[ICache.scala 27:22]
  reg  way0V_18; // @[ICache.scala 27:22]
  reg  way0V_19; // @[ICache.scala 27:22]
  reg  way0V_20; // @[ICache.scala 27:22]
  reg  way0V_21; // @[ICache.scala 27:22]
  reg  way0V_22; // @[ICache.scala 27:22]
  reg  way0V_23; // @[ICache.scala 27:22]
  reg  way0V_24; // @[ICache.scala 27:22]
  reg  way0V_25; // @[ICache.scala 27:22]
  reg  way0V_26; // @[ICache.scala 27:22]
  reg  way0V_27; // @[ICache.scala 27:22]
  reg  way0V_28; // @[ICache.scala 27:22]
  reg  way0V_29; // @[ICache.scala 27:22]
  reg  way0V_30; // @[ICache.scala 27:22]
  reg  way0V_31; // @[ICache.scala 27:22]
  reg  way0V_32; // @[ICache.scala 27:22]
  reg  way0V_33; // @[ICache.scala 27:22]
  reg  way0V_34; // @[ICache.scala 27:22]
  reg  way0V_35; // @[ICache.scala 27:22]
  reg  way0V_36; // @[ICache.scala 27:22]
  reg  way0V_37; // @[ICache.scala 27:22]
  reg  way0V_38; // @[ICache.scala 27:22]
  reg  way0V_39; // @[ICache.scala 27:22]
  reg  way0V_40; // @[ICache.scala 27:22]
  reg  way0V_41; // @[ICache.scala 27:22]
  reg  way0V_42; // @[ICache.scala 27:22]
  reg  way0V_43; // @[ICache.scala 27:22]
  reg  way0V_44; // @[ICache.scala 27:22]
  reg  way0V_45; // @[ICache.scala 27:22]
  reg  way0V_46; // @[ICache.scala 27:22]
  reg  way0V_47; // @[ICache.scala 27:22]
  reg  way0V_48; // @[ICache.scala 27:22]
  reg  way0V_49; // @[ICache.scala 27:22]
  reg  way0V_50; // @[ICache.scala 27:22]
  reg  way0V_51; // @[ICache.scala 27:22]
  reg  way0V_52; // @[ICache.scala 27:22]
  reg  way0V_53; // @[ICache.scala 27:22]
  reg  way0V_54; // @[ICache.scala 27:22]
  reg  way0V_55; // @[ICache.scala 27:22]
  reg  way0V_56; // @[ICache.scala 27:22]
  reg  way0V_57; // @[ICache.scala 27:22]
  reg  way0V_58; // @[ICache.scala 27:22]
  reg  way0V_59; // @[ICache.scala 27:22]
  reg  way0V_60; // @[ICache.scala 27:22]
  reg  way0V_61; // @[ICache.scala 27:22]
  reg  way0V_62; // @[ICache.scala 27:22]
  reg  way0V_63; // @[ICache.scala 27:22]
  reg  way0V_64; // @[ICache.scala 27:22]
  reg  way0V_65; // @[ICache.scala 27:22]
  reg  way0V_66; // @[ICache.scala 27:22]
  reg  way0V_67; // @[ICache.scala 27:22]
  reg  way0V_68; // @[ICache.scala 27:22]
  reg  way0V_69; // @[ICache.scala 27:22]
  reg  way0V_70; // @[ICache.scala 27:22]
  reg  way0V_71; // @[ICache.scala 27:22]
  reg  way0V_72; // @[ICache.scala 27:22]
  reg  way0V_73; // @[ICache.scala 27:22]
  reg  way0V_74; // @[ICache.scala 27:22]
  reg  way0V_75; // @[ICache.scala 27:22]
  reg  way0V_76; // @[ICache.scala 27:22]
  reg  way0V_77; // @[ICache.scala 27:22]
  reg  way0V_78; // @[ICache.scala 27:22]
  reg  way0V_79; // @[ICache.scala 27:22]
  reg  way0V_80; // @[ICache.scala 27:22]
  reg  way0V_81; // @[ICache.scala 27:22]
  reg  way0V_82; // @[ICache.scala 27:22]
  reg  way0V_83; // @[ICache.scala 27:22]
  reg  way0V_84; // @[ICache.scala 27:22]
  reg  way0V_85; // @[ICache.scala 27:22]
  reg  way0V_86; // @[ICache.scala 27:22]
  reg  way0V_87; // @[ICache.scala 27:22]
  reg  way0V_88; // @[ICache.scala 27:22]
  reg  way0V_89; // @[ICache.scala 27:22]
  reg  way0V_90; // @[ICache.scala 27:22]
  reg  way0V_91; // @[ICache.scala 27:22]
  reg  way0V_92; // @[ICache.scala 27:22]
  reg  way0V_93; // @[ICache.scala 27:22]
  reg  way0V_94; // @[ICache.scala 27:22]
  reg  way0V_95; // @[ICache.scala 27:22]
  reg  way0V_96; // @[ICache.scala 27:22]
  reg  way0V_97; // @[ICache.scala 27:22]
  reg  way0V_98; // @[ICache.scala 27:22]
  reg  way0V_99; // @[ICache.scala 27:22]
  reg  way0V_100; // @[ICache.scala 27:22]
  reg  way0V_101; // @[ICache.scala 27:22]
  reg  way0V_102; // @[ICache.scala 27:22]
  reg  way0V_103; // @[ICache.scala 27:22]
  reg  way0V_104; // @[ICache.scala 27:22]
  reg  way0V_105; // @[ICache.scala 27:22]
  reg  way0V_106; // @[ICache.scala 27:22]
  reg  way0V_107; // @[ICache.scala 27:22]
  reg  way0V_108; // @[ICache.scala 27:22]
  reg  way0V_109; // @[ICache.scala 27:22]
  reg  way0V_110; // @[ICache.scala 27:22]
  reg  way0V_111; // @[ICache.scala 27:22]
  reg  way0V_112; // @[ICache.scala 27:22]
  reg  way0V_113; // @[ICache.scala 27:22]
  reg  way0V_114; // @[ICache.scala 27:22]
  reg  way0V_115; // @[ICache.scala 27:22]
  reg  way0V_116; // @[ICache.scala 27:22]
  reg  way0V_117; // @[ICache.scala 27:22]
  reg  way0V_118; // @[ICache.scala 27:22]
  reg  way0V_119; // @[ICache.scala 27:22]
  reg  way0V_120; // @[ICache.scala 27:22]
  reg  way0V_121; // @[ICache.scala 27:22]
  reg  way0V_122; // @[ICache.scala 27:22]
  reg  way0V_123; // @[ICache.scala 27:22]
  reg  way0V_124; // @[ICache.scala 27:22]
  reg  way0V_125; // @[ICache.scala 27:22]
  reg  way0V_126; // @[ICache.scala 27:22]
  reg  way0V_127; // @[ICache.scala 27:22]
  reg [20:0] way0Tag_0; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_1; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_2; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_3; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_4; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_5; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_6; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_7; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_8; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_9; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_10; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_11; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_12; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_13; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_14; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_15; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_16; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_17; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_18; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_19; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_20; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_21; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_22; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_23; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_24; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_25; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_26; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_27; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_28; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_29; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_30; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_31; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_32; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_33; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_34; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_35; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_36; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_37; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_38; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_39; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_40; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_41; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_42; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_43; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_44; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_45; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_46; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_47; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_48; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_49; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_50; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_51; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_52; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_53; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_54; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_55; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_56; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_57; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_58; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_59; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_60; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_61; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_62; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_63; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_64; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_65; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_66; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_67; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_68; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_69; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_70; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_71; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_72; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_73; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_74; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_75; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_76; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_77; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_78; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_79; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_80; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_81; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_82; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_83; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_84; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_85; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_86; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_87; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_88; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_89; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_90; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_91; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_92; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_93; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_94; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_95; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_96; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_97; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_98; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_99; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_100; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_101; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_102; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_103; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_104; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_105; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_106; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_107; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_108; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_109; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_110; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_111; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_112; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_113; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_114; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_115; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_116; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_117; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_118; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_119; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_120; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_121; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_122; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_123; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_124; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_125; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_126; // @[ICache.scala 28:24]
  reg [20:0] way0Tag_127; // @[ICache.scala 28:24]
  reg  way0Age_0; // @[ICache.scala 30:24]
  reg  way0Age_1; // @[ICache.scala 30:24]
  reg  way0Age_2; // @[ICache.scala 30:24]
  reg  way0Age_3; // @[ICache.scala 30:24]
  reg  way0Age_4; // @[ICache.scala 30:24]
  reg  way0Age_5; // @[ICache.scala 30:24]
  reg  way0Age_6; // @[ICache.scala 30:24]
  reg  way0Age_7; // @[ICache.scala 30:24]
  reg  way0Age_8; // @[ICache.scala 30:24]
  reg  way0Age_9; // @[ICache.scala 30:24]
  reg  way0Age_10; // @[ICache.scala 30:24]
  reg  way0Age_11; // @[ICache.scala 30:24]
  reg  way0Age_12; // @[ICache.scala 30:24]
  reg  way0Age_13; // @[ICache.scala 30:24]
  reg  way0Age_14; // @[ICache.scala 30:24]
  reg  way0Age_15; // @[ICache.scala 30:24]
  reg  way0Age_16; // @[ICache.scala 30:24]
  reg  way0Age_17; // @[ICache.scala 30:24]
  reg  way0Age_18; // @[ICache.scala 30:24]
  reg  way0Age_19; // @[ICache.scala 30:24]
  reg  way0Age_20; // @[ICache.scala 30:24]
  reg  way0Age_21; // @[ICache.scala 30:24]
  reg  way0Age_22; // @[ICache.scala 30:24]
  reg  way0Age_23; // @[ICache.scala 30:24]
  reg  way0Age_24; // @[ICache.scala 30:24]
  reg  way0Age_25; // @[ICache.scala 30:24]
  reg  way0Age_26; // @[ICache.scala 30:24]
  reg  way0Age_27; // @[ICache.scala 30:24]
  reg  way0Age_28; // @[ICache.scala 30:24]
  reg  way0Age_29; // @[ICache.scala 30:24]
  reg  way0Age_30; // @[ICache.scala 30:24]
  reg  way0Age_31; // @[ICache.scala 30:24]
  reg  way0Age_32; // @[ICache.scala 30:24]
  reg  way0Age_33; // @[ICache.scala 30:24]
  reg  way0Age_34; // @[ICache.scala 30:24]
  reg  way0Age_35; // @[ICache.scala 30:24]
  reg  way0Age_36; // @[ICache.scala 30:24]
  reg  way0Age_37; // @[ICache.scala 30:24]
  reg  way0Age_38; // @[ICache.scala 30:24]
  reg  way0Age_39; // @[ICache.scala 30:24]
  reg  way0Age_40; // @[ICache.scala 30:24]
  reg  way0Age_41; // @[ICache.scala 30:24]
  reg  way0Age_42; // @[ICache.scala 30:24]
  reg  way0Age_43; // @[ICache.scala 30:24]
  reg  way0Age_44; // @[ICache.scala 30:24]
  reg  way0Age_45; // @[ICache.scala 30:24]
  reg  way0Age_46; // @[ICache.scala 30:24]
  reg  way0Age_47; // @[ICache.scala 30:24]
  reg  way0Age_48; // @[ICache.scala 30:24]
  reg  way0Age_49; // @[ICache.scala 30:24]
  reg  way0Age_50; // @[ICache.scala 30:24]
  reg  way0Age_51; // @[ICache.scala 30:24]
  reg  way0Age_52; // @[ICache.scala 30:24]
  reg  way0Age_53; // @[ICache.scala 30:24]
  reg  way0Age_54; // @[ICache.scala 30:24]
  reg  way0Age_55; // @[ICache.scala 30:24]
  reg  way0Age_56; // @[ICache.scala 30:24]
  reg  way0Age_57; // @[ICache.scala 30:24]
  reg  way0Age_58; // @[ICache.scala 30:24]
  reg  way0Age_59; // @[ICache.scala 30:24]
  reg  way0Age_60; // @[ICache.scala 30:24]
  reg  way0Age_61; // @[ICache.scala 30:24]
  reg  way0Age_62; // @[ICache.scala 30:24]
  reg  way0Age_63; // @[ICache.scala 30:24]
  reg  way0Age_64; // @[ICache.scala 30:24]
  reg  way0Age_65; // @[ICache.scala 30:24]
  reg  way0Age_66; // @[ICache.scala 30:24]
  reg  way0Age_67; // @[ICache.scala 30:24]
  reg  way0Age_68; // @[ICache.scala 30:24]
  reg  way0Age_69; // @[ICache.scala 30:24]
  reg  way0Age_70; // @[ICache.scala 30:24]
  reg  way0Age_71; // @[ICache.scala 30:24]
  reg  way0Age_72; // @[ICache.scala 30:24]
  reg  way0Age_73; // @[ICache.scala 30:24]
  reg  way0Age_74; // @[ICache.scala 30:24]
  reg  way0Age_75; // @[ICache.scala 30:24]
  reg  way0Age_76; // @[ICache.scala 30:24]
  reg  way0Age_77; // @[ICache.scala 30:24]
  reg  way0Age_78; // @[ICache.scala 30:24]
  reg  way0Age_79; // @[ICache.scala 30:24]
  reg  way0Age_80; // @[ICache.scala 30:24]
  reg  way0Age_81; // @[ICache.scala 30:24]
  reg  way0Age_82; // @[ICache.scala 30:24]
  reg  way0Age_83; // @[ICache.scala 30:24]
  reg  way0Age_84; // @[ICache.scala 30:24]
  reg  way0Age_85; // @[ICache.scala 30:24]
  reg  way0Age_86; // @[ICache.scala 30:24]
  reg  way0Age_87; // @[ICache.scala 30:24]
  reg  way0Age_88; // @[ICache.scala 30:24]
  reg  way0Age_89; // @[ICache.scala 30:24]
  reg  way0Age_90; // @[ICache.scala 30:24]
  reg  way0Age_91; // @[ICache.scala 30:24]
  reg  way0Age_92; // @[ICache.scala 30:24]
  reg  way0Age_93; // @[ICache.scala 30:24]
  reg  way0Age_94; // @[ICache.scala 30:24]
  reg  way0Age_95; // @[ICache.scala 30:24]
  reg  way0Age_96; // @[ICache.scala 30:24]
  reg  way0Age_97; // @[ICache.scala 30:24]
  reg  way0Age_98; // @[ICache.scala 30:24]
  reg  way0Age_99; // @[ICache.scala 30:24]
  reg  way0Age_100; // @[ICache.scala 30:24]
  reg  way0Age_101; // @[ICache.scala 30:24]
  reg  way0Age_102; // @[ICache.scala 30:24]
  reg  way0Age_103; // @[ICache.scala 30:24]
  reg  way0Age_104; // @[ICache.scala 30:24]
  reg  way0Age_105; // @[ICache.scala 30:24]
  reg  way0Age_106; // @[ICache.scala 30:24]
  reg  way0Age_107; // @[ICache.scala 30:24]
  reg  way0Age_108; // @[ICache.scala 30:24]
  reg  way0Age_109; // @[ICache.scala 30:24]
  reg  way0Age_110; // @[ICache.scala 30:24]
  reg  way0Age_111; // @[ICache.scala 30:24]
  reg  way0Age_112; // @[ICache.scala 30:24]
  reg  way0Age_113; // @[ICache.scala 30:24]
  reg  way0Age_114; // @[ICache.scala 30:24]
  reg  way0Age_115; // @[ICache.scala 30:24]
  reg  way0Age_116; // @[ICache.scala 30:24]
  reg  way0Age_117; // @[ICache.scala 30:24]
  reg  way0Age_118; // @[ICache.scala 30:24]
  reg  way0Age_119; // @[ICache.scala 30:24]
  reg  way0Age_120; // @[ICache.scala 30:24]
  reg  way0Age_121; // @[ICache.scala 30:24]
  reg  way0Age_122; // @[ICache.scala 30:24]
  reg  way0Age_123; // @[ICache.scala 30:24]
  reg  way0Age_124; // @[ICache.scala 30:24]
  reg  way0Age_125; // @[ICache.scala 30:24]
  reg  way0Age_126; // @[ICache.scala 30:24]
  reg  way0Age_127; // @[ICache.scala 30:24]
  reg  way1V_0; // @[ICache.scala 32:22]
  reg  way1V_1; // @[ICache.scala 32:22]
  reg  way1V_2; // @[ICache.scala 32:22]
  reg  way1V_3; // @[ICache.scala 32:22]
  reg  way1V_4; // @[ICache.scala 32:22]
  reg  way1V_5; // @[ICache.scala 32:22]
  reg  way1V_6; // @[ICache.scala 32:22]
  reg  way1V_7; // @[ICache.scala 32:22]
  reg  way1V_8; // @[ICache.scala 32:22]
  reg  way1V_9; // @[ICache.scala 32:22]
  reg  way1V_10; // @[ICache.scala 32:22]
  reg  way1V_11; // @[ICache.scala 32:22]
  reg  way1V_12; // @[ICache.scala 32:22]
  reg  way1V_13; // @[ICache.scala 32:22]
  reg  way1V_14; // @[ICache.scala 32:22]
  reg  way1V_15; // @[ICache.scala 32:22]
  reg  way1V_16; // @[ICache.scala 32:22]
  reg  way1V_17; // @[ICache.scala 32:22]
  reg  way1V_18; // @[ICache.scala 32:22]
  reg  way1V_19; // @[ICache.scala 32:22]
  reg  way1V_20; // @[ICache.scala 32:22]
  reg  way1V_21; // @[ICache.scala 32:22]
  reg  way1V_22; // @[ICache.scala 32:22]
  reg  way1V_23; // @[ICache.scala 32:22]
  reg  way1V_24; // @[ICache.scala 32:22]
  reg  way1V_25; // @[ICache.scala 32:22]
  reg  way1V_26; // @[ICache.scala 32:22]
  reg  way1V_27; // @[ICache.scala 32:22]
  reg  way1V_28; // @[ICache.scala 32:22]
  reg  way1V_29; // @[ICache.scala 32:22]
  reg  way1V_30; // @[ICache.scala 32:22]
  reg  way1V_31; // @[ICache.scala 32:22]
  reg  way1V_32; // @[ICache.scala 32:22]
  reg  way1V_33; // @[ICache.scala 32:22]
  reg  way1V_34; // @[ICache.scala 32:22]
  reg  way1V_35; // @[ICache.scala 32:22]
  reg  way1V_36; // @[ICache.scala 32:22]
  reg  way1V_37; // @[ICache.scala 32:22]
  reg  way1V_38; // @[ICache.scala 32:22]
  reg  way1V_39; // @[ICache.scala 32:22]
  reg  way1V_40; // @[ICache.scala 32:22]
  reg  way1V_41; // @[ICache.scala 32:22]
  reg  way1V_42; // @[ICache.scala 32:22]
  reg  way1V_43; // @[ICache.scala 32:22]
  reg  way1V_44; // @[ICache.scala 32:22]
  reg  way1V_45; // @[ICache.scala 32:22]
  reg  way1V_46; // @[ICache.scala 32:22]
  reg  way1V_47; // @[ICache.scala 32:22]
  reg  way1V_48; // @[ICache.scala 32:22]
  reg  way1V_49; // @[ICache.scala 32:22]
  reg  way1V_50; // @[ICache.scala 32:22]
  reg  way1V_51; // @[ICache.scala 32:22]
  reg  way1V_52; // @[ICache.scala 32:22]
  reg  way1V_53; // @[ICache.scala 32:22]
  reg  way1V_54; // @[ICache.scala 32:22]
  reg  way1V_55; // @[ICache.scala 32:22]
  reg  way1V_56; // @[ICache.scala 32:22]
  reg  way1V_57; // @[ICache.scala 32:22]
  reg  way1V_58; // @[ICache.scala 32:22]
  reg  way1V_59; // @[ICache.scala 32:22]
  reg  way1V_60; // @[ICache.scala 32:22]
  reg  way1V_61; // @[ICache.scala 32:22]
  reg  way1V_62; // @[ICache.scala 32:22]
  reg  way1V_63; // @[ICache.scala 32:22]
  reg  way1V_64; // @[ICache.scala 32:22]
  reg  way1V_65; // @[ICache.scala 32:22]
  reg  way1V_66; // @[ICache.scala 32:22]
  reg  way1V_67; // @[ICache.scala 32:22]
  reg  way1V_68; // @[ICache.scala 32:22]
  reg  way1V_69; // @[ICache.scala 32:22]
  reg  way1V_70; // @[ICache.scala 32:22]
  reg  way1V_71; // @[ICache.scala 32:22]
  reg  way1V_72; // @[ICache.scala 32:22]
  reg  way1V_73; // @[ICache.scala 32:22]
  reg  way1V_74; // @[ICache.scala 32:22]
  reg  way1V_75; // @[ICache.scala 32:22]
  reg  way1V_76; // @[ICache.scala 32:22]
  reg  way1V_77; // @[ICache.scala 32:22]
  reg  way1V_78; // @[ICache.scala 32:22]
  reg  way1V_79; // @[ICache.scala 32:22]
  reg  way1V_80; // @[ICache.scala 32:22]
  reg  way1V_81; // @[ICache.scala 32:22]
  reg  way1V_82; // @[ICache.scala 32:22]
  reg  way1V_83; // @[ICache.scala 32:22]
  reg  way1V_84; // @[ICache.scala 32:22]
  reg  way1V_85; // @[ICache.scala 32:22]
  reg  way1V_86; // @[ICache.scala 32:22]
  reg  way1V_87; // @[ICache.scala 32:22]
  reg  way1V_88; // @[ICache.scala 32:22]
  reg  way1V_89; // @[ICache.scala 32:22]
  reg  way1V_90; // @[ICache.scala 32:22]
  reg  way1V_91; // @[ICache.scala 32:22]
  reg  way1V_92; // @[ICache.scala 32:22]
  reg  way1V_93; // @[ICache.scala 32:22]
  reg  way1V_94; // @[ICache.scala 32:22]
  reg  way1V_95; // @[ICache.scala 32:22]
  reg  way1V_96; // @[ICache.scala 32:22]
  reg  way1V_97; // @[ICache.scala 32:22]
  reg  way1V_98; // @[ICache.scala 32:22]
  reg  way1V_99; // @[ICache.scala 32:22]
  reg  way1V_100; // @[ICache.scala 32:22]
  reg  way1V_101; // @[ICache.scala 32:22]
  reg  way1V_102; // @[ICache.scala 32:22]
  reg  way1V_103; // @[ICache.scala 32:22]
  reg  way1V_104; // @[ICache.scala 32:22]
  reg  way1V_105; // @[ICache.scala 32:22]
  reg  way1V_106; // @[ICache.scala 32:22]
  reg  way1V_107; // @[ICache.scala 32:22]
  reg  way1V_108; // @[ICache.scala 32:22]
  reg  way1V_109; // @[ICache.scala 32:22]
  reg  way1V_110; // @[ICache.scala 32:22]
  reg  way1V_111; // @[ICache.scala 32:22]
  reg  way1V_112; // @[ICache.scala 32:22]
  reg  way1V_113; // @[ICache.scala 32:22]
  reg  way1V_114; // @[ICache.scala 32:22]
  reg  way1V_115; // @[ICache.scala 32:22]
  reg  way1V_116; // @[ICache.scala 32:22]
  reg  way1V_117; // @[ICache.scala 32:22]
  reg  way1V_118; // @[ICache.scala 32:22]
  reg  way1V_119; // @[ICache.scala 32:22]
  reg  way1V_120; // @[ICache.scala 32:22]
  reg  way1V_121; // @[ICache.scala 32:22]
  reg  way1V_122; // @[ICache.scala 32:22]
  reg  way1V_123; // @[ICache.scala 32:22]
  reg  way1V_124; // @[ICache.scala 32:22]
  reg  way1V_125; // @[ICache.scala 32:22]
  reg  way1V_126; // @[ICache.scala 32:22]
  reg  way1V_127; // @[ICache.scala 32:22]
  reg [20:0] way1Tag_0; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_1; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_2; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_3; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_4; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_5; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_6; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_7; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_8; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_9; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_10; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_11; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_12; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_13; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_14; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_15; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_16; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_17; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_18; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_19; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_20; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_21; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_22; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_23; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_24; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_25; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_26; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_27; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_28; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_29; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_30; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_31; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_32; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_33; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_34; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_35; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_36; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_37; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_38; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_39; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_40; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_41; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_42; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_43; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_44; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_45; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_46; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_47; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_48; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_49; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_50; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_51; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_52; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_53; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_54; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_55; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_56; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_57; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_58; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_59; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_60; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_61; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_62; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_63; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_64; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_65; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_66; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_67; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_68; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_69; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_70; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_71; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_72; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_73; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_74; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_75; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_76; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_77; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_78; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_79; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_80; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_81; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_82; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_83; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_84; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_85; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_86; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_87; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_88; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_89; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_90; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_91; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_92; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_93; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_94; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_95; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_96; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_97; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_98; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_99; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_100; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_101; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_102; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_103; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_104; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_105; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_106; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_107; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_108; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_109; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_110; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_111; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_112; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_113; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_114; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_115; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_116; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_117; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_118; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_119; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_120; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_121; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_122; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_123; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_124; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_125; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_126; // @[ICache.scala 33:24]
  reg [20:0] way1Tag_127; // @[ICache.scala 33:24]
  reg  way1Age_0; // @[ICache.scala 35:24]
  reg  way1Age_1; // @[ICache.scala 35:24]
  reg  way1Age_2; // @[ICache.scala 35:24]
  reg  way1Age_3; // @[ICache.scala 35:24]
  reg  way1Age_4; // @[ICache.scala 35:24]
  reg  way1Age_5; // @[ICache.scala 35:24]
  reg  way1Age_6; // @[ICache.scala 35:24]
  reg  way1Age_7; // @[ICache.scala 35:24]
  reg  way1Age_8; // @[ICache.scala 35:24]
  reg  way1Age_9; // @[ICache.scala 35:24]
  reg  way1Age_10; // @[ICache.scala 35:24]
  reg  way1Age_11; // @[ICache.scala 35:24]
  reg  way1Age_12; // @[ICache.scala 35:24]
  reg  way1Age_13; // @[ICache.scala 35:24]
  reg  way1Age_14; // @[ICache.scala 35:24]
  reg  way1Age_15; // @[ICache.scala 35:24]
  reg  way1Age_16; // @[ICache.scala 35:24]
  reg  way1Age_17; // @[ICache.scala 35:24]
  reg  way1Age_18; // @[ICache.scala 35:24]
  reg  way1Age_19; // @[ICache.scala 35:24]
  reg  way1Age_20; // @[ICache.scala 35:24]
  reg  way1Age_21; // @[ICache.scala 35:24]
  reg  way1Age_22; // @[ICache.scala 35:24]
  reg  way1Age_23; // @[ICache.scala 35:24]
  reg  way1Age_24; // @[ICache.scala 35:24]
  reg  way1Age_25; // @[ICache.scala 35:24]
  reg  way1Age_26; // @[ICache.scala 35:24]
  reg  way1Age_27; // @[ICache.scala 35:24]
  reg  way1Age_28; // @[ICache.scala 35:24]
  reg  way1Age_29; // @[ICache.scala 35:24]
  reg  way1Age_30; // @[ICache.scala 35:24]
  reg  way1Age_31; // @[ICache.scala 35:24]
  reg  way1Age_32; // @[ICache.scala 35:24]
  reg  way1Age_33; // @[ICache.scala 35:24]
  reg  way1Age_34; // @[ICache.scala 35:24]
  reg  way1Age_35; // @[ICache.scala 35:24]
  reg  way1Age_36; // @[ICache.scala 35:24]
  reg  way1Age_37; // @[ICache.scala 35:24]
  reg  way1Age_38; // @[ICache.scala 35:24]
  reg  way1Age_39; // @[ICache.scala 35:24]
  reg  way1Age_40; // @[ICache.scala 35:24]
  reg  way1Age_41; // @[ICache.scala 35:24]
  reg  way1Age_42; // @[ICache.scala 35:24]
  reg  way1Age_43; // @[ICache.scala 35:24]
  reg  way1Age_44; // @[ICache.scala 35:24]
  reg  way1Age_45; // @[ICache.scala 35:24]
  reg  way1Age_46; // @[ICache.scala 35:24]
  reg  way1Age_47; // @[ICache.scala 35:24]
  reg  way1Age_48; // @[ICache.scala 35:24]
  reg  way1Age_49; // @[ICache.scala 35:24]
  reg  way1Age_50; // @[ICache.scala 35:24]
  reg  way1Age_51; // @[ICache.scala 35:24]
  reg  way1Age_52; // @[ICache.scala 35:24]
  reg  way1Age_53; // @[ICache.scala 35:24]
  reg  way1Age_54; // @[ICache.scala 35:24]
  reg  way1Age_55; // @[ICache.scala 35:24]
  reg  way1Age_56; // @[ICache.scala 35:24]
  reg  way1Age_57; // @[ICache.scala 35:24]
  reg  way1Age_58; // @[ICache.scala 35:24]
  reg  way1Age_59; // @[ICache.scala 35:24]
  reg  way1Age_60; // @[ICache.scala 35:24]
  reg  way1Age_61; // @[ICache.scala 35:24]
  reg  way1Age_62; // @[ICache.scala 35:24]
  reg  way1Age_63; // @[ICache.scala 35:24]
  reg  way1Age_64; // @[ICache.scala 35:24]
  reg  way1Age_65; // @[ICache.scala 35:24]
  reg  way1Age_66; // @[ICache.scala 35:24]
  reg  way1Age_67; // @[ICache.scala 35:24]
  reg  way1Age_68; // @[ICache.scala 35:24]
  reg  way1Age_69; // @[ICache.scala 35:24]
  reg  way1Age_70; // @[ICache.scala 35:24]
  reg  way1Age_71; // @[ICache.scala 35:24]
  reg  way1Age_72; // @[ICache.scala 35:24]
  reg  way1Age_73; // @[ICache.scala 35:24]
  reg  way1Age_74; // @[ICache.scala 35:24]
  reg  way1Age_75; // @[ICache.scala 35:24]
  reg  way1Age_76; // @[ICache.scala 35:24]
  reg  way1Age_77; // @[ICache.scala 35:24]
  reg  way1Age_78; // @[ICache.scala 35:24]
  reg  way1Age_79; // @[ICache.scala 35:24]
  reg  way1Age_80; // @[ICache.scala 35:24]
  reg  way1Age_81; // @[ICache.scala 35:24]
  reg  way1Age_82; // @[ICache.scala 35:24]
  reg  way1Age_83; // @[ICache.scala 35:24]
  reg  way1Age_84; // @[ICache.scala 35:24]
  reg  way1Age_85; // @[ICache.scala 35:24]
  reg  way1Age_86; // @[ICache.scala 35:24]
  reg  way1Age_87; // @[ICache.scala 35:24]
  reg  way1Age_88; // @[ICache.scala 35:24]
  reg  way1Age_89; // @[ICache.scala 35:24]
  reg  way1Age_90; // @[ICache.scala 35:24]
  reg  way1Age_91; // @[ICache.scala 35:24]
  reg  way1Age_92; // @[ICache.scala 35:24]
  reg  way1Age_93; // @[ICache.scala 35:24]
  reg  way1Age_94; // @[ICache.scala 35:24]
  reg  way1Age_95; // @[ICache.scala 35:24]
  reg  way1Age_96; // @[ICache.scala 35:24]
  reg  way1Age_97; // @[ICache.scala 35:24]
  reg  way1Age_98; // @[ICache.scala 35:24]
  reg  way1Age_99; // @[ICache.scala 35:24]
  reg  way1Age_100; // @[ICache.scala 35:24]
  reg  way1Age_101; // @[ICache.scala 35:24]
  reg  way1Age_102; // @[ICache.scala 35:24]
  reg  way1Age_103; // @[ICache.scala 35:24]
  reg  way1Age_104; // @[ICache.scala 35:24]
  reg  way1Age_105; // @[ICache.scala 35:24]
  reg  way1Age_106; // @[ICache.scala 35:24]
  reg  way1Age_107; // @[ICache.scala 35:24]
  reg  way1Age_108; // @[ICache.scala 35:24]
  reg  way1Age_109; // @[ICache.scala 35:24]
  reg  way1Age_110; // @[ICache.scala 35:24]
  reg  way1Age_111; // @[ICache.scala 35:24]
  reg  way1Age_112; // @[ICache.scala 35:24]
  reg  way1Age_113; // @[ICache.scala 35:24]
  reg  way1Age_114; // @[ICache.scala 35:24]
  reg  way1Age_115; // @[ICache.scala 35:24]
  reg  way1Age_116; // @[ICache.scala 35:24]
  reg  way1Age_117; // @[ICache.scala 35:24]
  reg  way1Age_118; // @[ICache.scala 35:24]
  reg  way1Age_119; // @[ICache.scala 35:24]
  reg  way1Age_120; // @[ICache.scala 35:24]
  reg  way1Age_121; // @[ICache.scala 35:24]
  reg  way1Age_122; // @[ICache.scala 35:24]
  reg  way1Age_123; // @[ICache.scala 35:24]
  reg  way1Age_124; // @[ICache.scala 35:24]
  reg  way1Age_125; // @[ICache.scala 35:24]
  reg  way1Age_126; // @[ICache.scala 35:24]
  reg  way1Age_127; // @[ICache.scala 35:24]
  reg [1:0] state; // @[ICache.scala 38:22]
  wire [20:0] reqTag = io_imem_inst_addr[31:11]; // @[ICache.scala 42:25]
  wire [6:0] reqIndex = io_imem_inst_addr[10:4]; // @[ICache.scala 43:27]
  wire [3:0] reqOff = io_imem_inst_addr[3:0]; // @[ICache.scala 44:25]
  wire [20:0] _GEN_1 = 7'h1 == reqIndex ? way0Tag_1 : way0Tag_0; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_2 = 7'h2 == reqIndex ? way0Tag_2 : _GEN_1; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_3 = 7'h3 == reqIndex ? way0Tag_3 : _GEN_2; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_4 = 7'h4 == reqIndex ? way0Tag_4 : _GEN_3; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_5 = 7'h5 == reqIndex ? way0Tag_5 : _GEN_4; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_6 = 7'h6 == reqIndex ? way0Tag_6 : _GEN_5; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_7 = 7'h7 == reqIndex ? way0Tag_7 : _GEN_6; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_8 = 7'h8 == reqIndex ? way0Tag_8 : _GEN_7; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_9 = 7'h9 == reqIndex ? way0Tag_9 : _GEN_8; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_10 = 7'ha == reqIndex ? way0Tag_10 : _GEN_9; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_11 = 7'hb == reqIndex ? way0Tag_11 : _GEN_10; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_12 = 7'hc == reqIndex ? way0Tag_12 : _GEN_11; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_13 = 7'hd == reqIndex ? way0Tag_13 : _GEN_12; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_14 = 7'he == reqIndex ? way0Tag_14 : _GEN_13; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_15 = 7'hf == reqIndex ? way0Tag_15 : _GEN_14; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_16 = 7'h10 == reqIndex ? way0Tag_16 : _GEN_15; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_17 = 7'h11 == reqIndex ? way0Tag_17 : _GEN_16; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_18 = 7'h12 == reqIndex ? way0Tag_18 : _GEN_17; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_19 = 7'h13 == reqIndex ? way0Tag_19 : _GEN_18; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_20 = 7'h14 == reqIndex ? way0Tag_20 : _GEN_19; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_21 = 7'h15 == reqIndex ? way0Tag_21 : _GEN_20; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_22 = 7'h16 == reqIndex ? way0Tag_22 : _GEN_21; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_23 = 7'h17 == reqIndex ? way0Tag_23 : _GEN_22; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_24 = 7'h18 == reqIndex ? way0Tag_24 : _GEN_23; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_25 = 7'h19 == reqIndex ? way0Tag_25 : _GEN_24; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_26 = 7'h1a == reqIndex ? way0Tag_26 : _GEN_25; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_27 = 7'h1b == reqIndex ? way0Tag_27 : _GEN_26; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_28 = 7'h1c == reqIndex ? way0Tag_28 : _GEN_27; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_29 = 7'h1d == reqIndex ? way0Tag_29 : _GEN_28; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_30 = 7'h1e == reqIndex ? way0Tag_30 : _GEN_29; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_31 = 7'h1f == reqIndex ? way0Tag_31 : _GEN_30; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_32 = 7'h20 == reqIndex ? way0Tag_32 : _GEN_31; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_33 = 7'h21 == reqIndex ? way0Tag_33 : _GEN_32; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_34 = 7'h22 == reqIndex ? way0Tag_34 : _GEN_33; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_35 = 7'h23 == reqIndex ? way0Tag_35 : _GEN_34; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_36 = 7'h24 == reqIndex ? way0Tag_36 : _GEN_35; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_37 = 7'h25 == reqIndex ? way0Tag_37 : _GEN_36; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_38 = 7'h26 == reqIndex ? way0Tag_38 : _GEN_37; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_39 = 7'h27 == reqIndex ? way0Tag_39 : _GEN_38; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_40 = 7'h28 == reqIndex ? way0Tag_40 : _GEN_39; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_41 = 7'h29 == reqIndex ? way0Tag_41 : _GEN_40; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_42 = 7'h2a == reqIndex ? way0Tag_42 : _GEN_41; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_43 = 7'h2b == reqIndex ? way0Tag_43 : _GEN_42; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_44 = 7'h2c == reqIndex ? way0Tag_44 : _GEN_43; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_45 = 7'h2d == reqIndex ? way0Tag_45 : _GEN_44; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_46 = 7'h2e == reqIndex ? way0Tag_46 : _GEN_45; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_47 = 7'h2f == reqIndex ? way0Tag_47 : _GEN_46; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_48 = 7'h30 == reqIndex ? way0Tag_48 : _GEN_47; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_49 = 7'h31 == reqIndex ? way0Tag_49 : _GEN_48; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_50 = 7'h32 == reqIndex ? way0Tag_50 : _GEN_49; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_51 = 7'h33 == reqIndex ? way0Tag_51 : _GEN_50; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_52 = 7'h34 == reqIndex ? way0Tag_52 : _GEN_51; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_53 = 7'h35 == reqIndex ? way0Tag_53 : _GEN_52; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_54 = 7'h36 == reqIndex ? way0Tag_54 : _GEN_53; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_55 = 7'h37 == reqIndex ? way0Tag_55 : _GEN_54; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_56 = 7'h38 == reqIndex ? way0Tag_56 : _GEN_55; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_57 = 7'h39 == reqIndex ? way0Tag_57 : _GEN_56; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_58 = 7'h3a == reqIndex ? way0Tag_58 : _GEN_57; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_59 = 7'h3b == reqIndex ? way0Tag_59 : _GEN_58; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_60 = 7'h3c == reqIndex ? way0Tag_60 : _GEN_59; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_61 = 7'h3d == reqIndex ? way0Tag_61 : _GEN_60; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_62 = 7'h3e == reqIndex ? way0Tag_62 : _GEN_61; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_63 = 7'h3f == reqIndex ? way0Tag_63 : _GEN_62; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_64 = 7'h40 == reqIndex ? way0Tag_64 : _GEN_63; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_65 = 7'h41 == reqIndex ? way0Tag_65 : _GEN_64; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_66 = 7'h42 == reqIndex ? way0Tag_66 : _GEN_65; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_67 = 7'h43 == reqIndex ? way0Tag_67 : _GEN_66; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_68 = 7'h44 == reqIndex ? way0Tag_68 : _GEN_67; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_69 = 7'h45 == reqIndex ? way0Tag_69 : _GEN_68; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_70 = 7'h46 == reqIndex ? way0Tag_70 : _GEN_69; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_71 = 7'h47 == reqIndex ? way0Tag_71 : _GEN_70; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_72 = 7'h48 == reqIndex ? way0Tag_72 : _GEN_71; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_73 = 7'h49 == reqIndex ? way0Tag_73 : _GEN_72; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_74 = 7'h4a == reqIndex ? way0Tag_74 : _GEN_73; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_75 = 7'h4b == reqIndex ? way0Tag_75 : _GEN_74; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_76 = 7'h4c == reqIndex ? way0Tag_76 : _GEN_75; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_77 = 7'h4d == reqIndex ? way0Tag_77 : _GEN_76; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_78 = 7'h4e == reqIndex ? way0Tag_78 : _GEN_77; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_79 = 7'h4f == reqIndex ? way0Tag_79 : _GEN_78; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_80 = 7'h50 == reqIndex ? way0Tag_80 : _GEN_79; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_81 = 7'h51 == reqIndex ? way0Tag_81 : _GEN_80; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_82 = 7'h52 == reqIndex ? way0Tag_82 : _GEN_81; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_83 = 7'h53 == reqIndex ? way0Tag_83 : _GEN_82; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_84 = 7'h54 == reqIndex ? way0Tag_84 : _GEN_83; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_85 = 7'h55 == reqIndex ? way0Tag_85 : _GEN_84; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_86 = 7'h56 == reqIndex ? way0Tag_86 : _GEN_85; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_87 = 7'h57 == reqIndex ? way0Tag_87 : _GEN_86; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_88 = 7'h58 == reqIndex ? way0Tag_88 : _GEN_87; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_89 = 7'h59 == reqIndex ? way0Tag_89 : _GEN_88; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_90 = 7'h5a == reqIndex ? way0Tag_90 : _GEN_89; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_91 = 7'h5b == reqIndex ? way0Tag_91 : _GEN_90; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_92 = 7'h5c == reqIndex ? way0Tag_92 : _GEN_91; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_93 = 7'h5d == reqIndex ? way0Tag_93 : _GEN_92; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_94 = 7'h5e == reqIndex ? way0Tag_94 : _GEN_93; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_95 = 7'h5f == reqIndex ? way0Tag_95 : _GEN_94; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_96 = 7'h60 == reqIndex ? way0Tag_96 : _GEN_95; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_97 = 7'h61 == reqIndex ? way0Tag_97 : _GEN_96; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_98 = 7'h62 == reqIndex ? way0Tag_98 : _GEN_97; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_99 = 7'h63 == reqIndex ? way0Tag_99 : _GEN_98; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_100 = 7'h64 == reqIndex ? way0Tag_100 : _GEN_99; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_101 = 7'h65 == reqIndex ? way0Tag_101 : _GEN_100; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_102 = 7'h66 == reqIndex ? way0Tag_102 : _GEN_101; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_103 = 7'h67 == reqIndex ? way0Tag_103 : _GEN_102; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_104 = 7'h68 == reqIndex ? way0Tag_104 : _GEN_103; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_105 = 7'h69 == reqIndex ? way0Tag_105 : _GEN_104; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_106 = 7'h6a == reqIndex ? way0Tag_106 : _GEN_105; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_107 = 7'h6b == reqIndex ? way0Tag_107 : _GEN_106; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_108 = 7'h6c == reqIndex ? way0Tag_108 : _GEN_107; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_109 = 7'h6d == reqIndex ? way0Tag_109 : _GEN_108; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_110 = 7'h6e == reqIndex ? way0Tag_110 : _GEN_109; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_111 = 7'h6f == reqIndex ? way0Tag_111 : _GEN_110; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_112 = 7'h70 == reqIndex ? way0Tag_112 : _GEN_111; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_113 = 7'h71 == reqIndex ? way0Tag_113 : _GEN_112; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_114 = 7'h72 == reqIndex ? way0Tag_114 : _GEN_113; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_115 = 7'h73 == reqIndex ? way0Tag_115 : _GEN_114; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_116 = 7'h74 == reqIndex ? way0Tag_116 : _GEN_115; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_117 = 7'h75 == reqIndex ? way0Tag_117 : _GEN_116; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_118 = 7'h76 == reqIndex ? way0Tag_118 : _GEN_117; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_119 = 7'h77 == reqIndex ? way0Tag_119 : _GEN_118; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_120 = 7'h78 == reqIndex ? way0Tag_120 : _GEN_119; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_121 = 7'h79 == reqIndex ? way0Tag_121 : _GEN_120; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_122 = 7'h7a == reqIndex ? way0Tag_122 : _GEN_121; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_123 = 7'h7b == reqIndex ? way0Tag_123 : _GEN_122; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_124 = 7'h7c == reqIndex ? way0Tag_124 : _GEN_123; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_125 = 7'h7d == reqIndex ? way0Tag_125 : _GEN_124; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_126 = 7'h7e == reqIndex ? way0Tag_126 : _GEN_125; // @[ICache.scala 48:{55,55}]
  wire [20:0] _GEN_127 = 7'h7f == reqIndex ? way0Tag_127 : _GEN_126; // @[ICache.scala 48:{55,55}]
  wire  _GEN_129 = 7'h1 == reqIndex ? way0V_1 : way0V_0; // @[ICache.scala 48:{33,33}]
  wire  _GEN_130 = 7'h2 == reqIndex ? way0V_2 : _GEN_129; // @[ICache.scala 48:{33,33}]
  wire  _GEN_131 = 7'h3 == reqIndex ? way0V_3 : _GEN_130; // @[ICache.scala 48:{33,33}]
  wire  _GEN_132 = 7'h4 == reqIndex ? way0V_4 : _GEN_131; // @[ICache.scala 48:{33,33}]
  wire  _GEN_133 = 7'h5 == reqIndex ? way0V_5 : _GEN_132; // @[ICache.scala 48:{33,33}]
  wire  _GEN_134 = 7'h6 == reqIndex ? way0V_6 : _GEN_133; // @[ICache.scala 48:{33,33}]
  wire  _GEN_135 = 7'h7 == reqIndex ? way0V_7 : _GEN_134; // @[ICache.scala 48:{33,33}]
  wire  _GEN_136 = 7'h8 == reqIndex ? way0V_8 : _GEN_135; // @[ICache.scala 48:{33,33}]
  wire  _GEN_137 = 7'h9 == reqIndex ? way0V_9 : _GEN_136; // @[ICache.scala 48:{33,33}]
  wire  _GEN_138 = 7'ha == reqIndex ? way0V_10 : _GEN_137; // @[ICache.scala 48:{33,33}]
  wire  _GEN_139 = 7'hb == reqIndex ? way0V_11 : _GEN_138; // @[ICache.scala 48:{33,33}]
  wire  _GEN_140 = 7'hc == reqIndex ? way0V_12 : _GEN_139; // @[ICache.scala 48:{33,33}]
  wire  _GEN_141 = 7'hd == reqIndex ? way0V_13 : _GEN_140; // @[ICache.scala 48:{33,33}]
  wire  _GEN_142 = 7'he == reqIndex ? way0V_14 : _GEN_141; // @[ICache.scala 48:{33,33}]
  wire  _GEN_143 = 7'hf == reqIndex ? way0V_15 : _GEN_142; // @[ICache.scala 48:{33,33}]
  wire  _GEN_144 = 7'h10 == reqIndex ? way0V_16 : _GEN_143; // @[ICache.scala 48:{33,33}]
  wire  _GEN_145 = 7'h11 == reqIndex ? way0V_17 : _GEN_144; // @[ICache.scala 48:{33,33}]
  wire  _GEN_146 = 7'h12 == reqIndex ? way0V_18 : _GEN_145; // @[ICache.scala 48:{33,33}]
  wire  _GEN_147 = 7'h13 == reqIndex ? way0V_19 : _GEN_146; // @[ICache.scala 48:{33,33}]
  wire  _GEN_148 = 7'h14 == reqIndex ? way0V_20 : _GEN_147; // @[ICache.scala 48:{33,33}]
  wire  _GEN_149 = 7'h15 == reqIndex ? way0V_21 : _GEN_148; // @[ICache.scala 48:{33,33}]
  wire  _GEN_150 = 7'h16 == reqIndex ? way0V_22 : _GEN_149; // @[ICache.scala 48:{33,33}]
  wire  _GEN_151 = 7'h17 == reqIndex ? way0V_23 : _GEN_150; // @[ICache.scala 48:{33,33}]
  wire  _GEN_152 = 7'h18 == reqIndex ? way0V_24 : _GEN_151; // @[ICache.scala 48:{33,33}]
  wire  _GEN_153 = 7'h19 == reqIndex ? way0V_25 : _GEN_152; // @[ICache.scala 48:{33,33}]
  wire  _GEN_154 = 7'h1a == reqIndex ? way0V_26 : _GEN_153; // @[ICache.scala 48:{33,33}]
  wire  _GEN_155 = 7'h1b == reqIndex ? way0V_27 : _GEN_154; // @[ICache.scala 48:{33,33}]
  wire  _GEN_156 = 7'h1c == reqIndex ? way0V_28 : _GEN_155; // @[ICache.scala 48:{33,33}]
  wire  _GEN_157 = 7'h1d == reqIndex ? way0V_29 : _GEN_156; // @[ICache.scala 48:{33,33}]
  wire  _GEN_158 = 7'h1e == reqIndex ? way0V_30 : _GEN_157; // @[ICache.scala 48:{33,33}]
  wire  _GEN_159 = 7'h1f == reqIndex ? way0V_31 : _GEN_158; // @[ICache.scala 48:{33,33}]
  wire  _GEN_160 = 7'h20 == reqIndex ? way0V_32 : _GEN_159; // @[ICache.scala 48:{33,33}]
  wire  _GEN_161 = 7'h21 == reqIndex ? way0V_33 : _GEN_160; // @[ICache.scala 48:{33,33}]
  wire  _GEN_162 = 7'h22 == reqIndex ? way0V_34 : _GEN_161; // @[ICache.scala 48:{33,33}]
  wire  _GEN_163 = 7'h23 == reqIndex ? way0V_35 : _GEN_162; // @[ICache.scala 48:{33,33}]
  wire  _GEN_164 = 7'h24 == reqIndex ? way0V_36 : _GEN_163; // @[ICache.scala 48:{33,33}]
  wire  _GEN_165 = 7'h25 == reqIndex ? way0V_37 : _GEN_164; // @[ICache.scala 48:{33,33}]
  wire  _GEN_166 = 7'h26 == reqIndex ? way0V_38 : _GEN_165; // @[ICache.scala 48:{33,33}]
  wire  _GEN_167 = 7'h27 == reqIndex ? way0V_39 : _GEN_166; // @[ICache.scala 48:{33,33}]
  wire  _GEN_168 = 7'h28 == reqIndex ? way0V_40 : _GEN_167; // @[ICache.scala 48:{33,33}]
  wire  _GEN_169 = 7'h29 == reqIndex ? way0V_41 : _GEN_168; // @[ICache.scala 48:{33,33}]
  wire  _GEN_170 = 7'h2a == reqIndex ? way0V_42 : _GEN_169; // @[ICache.scala 48:{33,33}]
  wire  _GEN_171 = 7'h2b == reqIndex ? way0V_43 : _GEN_170; // @[ICache.scala 48:{33,33}]
  wire  _GEN_172 = 7'h2c == reqIndex ? way0V_44 : _GEN_171; // @[ICache.scala 48:{33,33}]
  wire  _GEN_173 = 7'h2d == reqIndex ? way0V_45 : _GEN_172; // @[ICache.scala 48:{33,33}]
  wire  _GEN_174 = 7'h2e == reqIndex ? way0V_46 : _GEN_173; // @[ICache.scala 48:{33,33}]
  wire  _GEN_175 = 7'h2f == reqIndex ? way0V_47 : _GEN_174; // @[ICache.scala 48:{33,33}]
  wire  _GEN_176 = 7'h30 == reqIndex ? way0V_48 : _GEN_175; // @[ICache.scala 48:{33,33}]
  wire  _GEN_177 = 7'h31 == reqIndex ? way0V_49 : _GEN_176; // @[ICache.scala 48:{33,33}]
  wire  _GEN_178 = 7'h32 == reqIndex ? way0V_50 : _GEN_177; // @[ICache.scala 48:{33,33}]
  wire  _GEN_179 = 7'h33 == reqIndex ? way0V_51 : _GEN_178; // @[ICache.scala 48:{33,33}]
  wire  _GEN_180 = 7'h34 == reqIndex ? way0V_52 : _GEN_179; // @[ICache.scala 48:{33,33}]
  wire  _GEN_181 = 7'h35 == reqIndex ? way0V_53 : _GEN_180; // @[ICache.scala 48:{33,33}]
  wire  _GEN_182 = 7'h36 == reqIndex ? way0V_54 : _GEN_181; // @[ICache.scala 48:{33,33}]
  wire  _GEN_183 = 7'h37 == reqIndex ? way0V_55 : _GEN_182; // @[ICache.scala 48:{33,33}]
  wire  _GEN_184 = 7'h38 == reqIndex ? way0V_56 : _GEN_183; // @[ICache.scala 48:{33,33}]
  wire  _GEN_185 = 7'h39 == reqIndex ? way0V_57 : _GEN_184; // @[ICache.scala 48:{33,33}]
  wire  _GEN_186 = 7'h3a == reqIndex ? way0V_58 : _GEN_185; // @[ICache.scala 48:{33,33}]
  wire  _GEN_187 = 7'h3b == reqIndex ? way0V_59 : _GEN_186; // @[ICache.scala 48:{33,33}]
  wire  _GEN_188 = 7'h3c == reqIndex ? way0V_60 : _GEN_187; // @[ICache.scala 48:{33,33}]
  wire  _GEN_189 = 7'h3d == reqIndex ? way0V_61 : _GEN_188; // @[ICache.scala 48:{33,33}]
  wire  _GEN_190 = 7'h3e == reqIndex ? way0V_62 : _GEN_189; // @[ICache.scala 48:{33,33}]
  wire  _GEN_191 = 7'h3f == reqIndex ? way0V_63 : _GEN_190; // @[ICache.scala 48:{33,33}]
  wire  _GEN_192 = 7'h40 == reqIndex ? way0V_64 : _GEN_191; // @[ICache.scala 48:{33,33}]
  wire  _GEN_193 = 7'h41 == reqIndex ? way0V_65 : _GEN_192; // @[ICache.scala 48:{33,33}]
  wire  _GEN_194 = 7'h42 == reqIndex ? way0V_66 : _GEN_193; // @[ICache.scala 48:{33,33}]
  wire  _GEN_195 = 7'h43 == reqIndex ? way0V_67 : _GEN_194; // @[ICache.scala 48:{33,33}]
  wire  _GEN_196 = 7'h44 == reqIndex ? way0V_68 : _GEN_195; // @[ICache.scala 48:{33,33}]
  wire  _GEN_197 = 7'h45 == reqIndex ? way0V_69 : _GEN_196; // @[ICache.scala 48:{33,33}]
  wire  _GEN_198 = 7'h46 == reqIndex ? way0V_70 : _GEN_197; // @[ICache.scala 48:{33,33}]
  wire  _GEN_199 = 7'h47 == reqIndex ? way0V_71 : _GEN_198; // @[ICache.scala 48:{33,33}]
  wire  _GEN_200 = 7'h48 == reqIndex ? way0V_72 : _GEN_199; // @[ICache.scala 48:{33,33}]
  wire  _GEN_201 = 7'h49 == reqIndex ? way0V_73 : _GEN_200; // @[ICache.scala 48:{33,33}]
  wire  _GEN_202 = 7'h4a == reqIndex ? way0V_74 : _GEN_201; // @[ICache.scala 48:{33,33}]
  wire  _GEN_203 = 7'h4b == reqIndex ? way0V_75 : _GEN_202; // @[ICache.scala 48:{33,33}]
  wire  _GEN_204 = 7'h4c == reqIndex ? way0V_76 : _GEN_203; // @[ICache.scala 48:{33,33}]
  wire  _GEN_205 = 7'h4d == reqIndex ? way0V_77 : _GEN_204; // @[ICache.scala 48:{33,33}]
  wire  _GEN_206 = 7'h4e == reqIndex ? way0V_78 : _GEN_205; // @[ICache.scala 48:{33,33}]
  wire  _GEN_207 = 7'h4f == reqIndex ? way0V_79 : _GEN_206; // @[ICache.scala 48:{33,33}]
  wire  _GEN_208 = 7'h50 == reqIndex ? way0V_80 : _GEN_207; // @[ICache.scala 48:{33,33}]
  wire  _GEN_209 = 7'h51 == reqIndex ? way0V_81 : _GEN_208; // @[ICache.scala 48:{33,33}]
  wire  _GEN_210 = 7'h52 == reqIndex ? way0V_82 : _GEN_209; // @[ICache.scala 48:{33,33}]
  wire  _GEN_211 = 7'h53 == reqIndex ? way0V_83 : _GEN_210; // @[ICache.scala 48:{33,33}]
  wire  _GEN_212 = 7'h54 == reqIndex ? way0V_84 : _GEN_211; // @[ICache.scala 48:{33,33}]
  wire  _GEN_213 = 7'h55 == reqIndex ? way0V_85 : _GEN_212; // @[ICache.scala 48:{33,33}]
  wire  _GEN_214 = 7'h56 == reqIndex ? way0V_86 : _GEN_213; // @[ICache.scala 48:{33,33}]
  wire  _GEN_215 = 7'h57 == reqIndex ? way0V_87 : _GEN_214; // @[ICache.scala 48:{33,33}]
  wire  _GEN_216 = 7'h58 == reqIndex ? way0V_88 : _GEN_215; // @[ICache.scala 48:{33,33}]
  wire  _GEN_217 = 7'h59 == reqIndex ? way0V_89 : _GEN_216; // @[ICache.scala 48:{33,33}]
  wire  _GEN_218 = 7'h5a == reqIndex ? way0V_90 : _GEN_217; // @[ICache.scala 48:{33,33}]
  wire  _GEN_219 = 7'h5b == reqIndex ? way0V_91 : _GEN_218; // @[ICache.scala 48:{33,33}]
  wire  _GEN_220 = 7'h5c == reqIndex ? way0V_92 : _GEN_219; // @[ICache.scala 48:{33,33}]
  wire  _GEN_221 = 7'h5d == reqIndex ? way0V_93 : _GEN_220; // @[ICache.scala 48:{33,33}]
  wire  _GEN_222 = 7'h5e == reqIndex ? way0V_94 : _GEN_221; // @[ICache.scala 48:{33,33}]
  wire  _GEN_223 = 7'h5f == reqIndex ? way0V_95 : _GEN_222; // @[ICache.scala 48:{33,33}]
  wire  _GEN_224 = 7'h60 == reqIndex ? way0V_96 : _GEN_223; // @[ICache.scala 48:{33,33}]
  wire  _GEN_225 = 7'h61 == reqIndex ? way0V_97 : _GEN_224; // @[ICache.scala 48:{33,33}]
  wire  _GEN_226 = 7'h62 == reqIndex ? way0V_98 : _GEN_225; // @[ICache.scala 48:{33,33}]
  wire  _GEN_227 = 7'h63 == reqIndex ? way0V_99 : _GEN_226; // @[ICache.scala 48:{33,33}]
  wire  _GEN_228 = 7'h64 == reqIndex ? way0V_100 : _GEN_227; // @[ICache.scala 48:{33,33}]
  wire  _GEN_229 = 7'h65 == reqIndex ? way0V_101 : _GEN_228; // @[ICache.scala 48:{33,33}]
  wire  _GEN_230 = 7'h66 == reqIndex ? way0V_102 : _GEN_229; // @[ICache.scala 48:{33,33}]
  wire  _GEN_231 = 7'h67 == reqIndex ? way0V_103 : _GEN_230; // @[ICache.scala 48:{33,33}]
  wire  _GEN_232 = 7'h68 == reqIndex ? way0V_104 : _GEN_231; // @[ICache.scala 48:{33,33}]
  wire  _GEN_233 = 7'h69 == reqIndex ? way0V_105 : _GEN_232; // @[ICache.scala 48:{33,33}]
  wire  _GEN_234 = 7'h6a == reqIndex ? way0V_106 : _GEN_233; // @[ICache.scala 48:{33,33}]
  wire  _GEN_235 = 7'h6b == reqIndex ? way0V_107 : _GEN_234; // @[ICache.scala 48:{33,33}]
  wire  _GEN_236 = 7'h6c == reqIndex ? way0V_108 : _GEN_235; // @[ICache.scala 48:{33,33}]
  wire  _GEN_237 = 7'h6d == reqIndex ? way0V_109 : _GEN_236; // @[ICache.scala 48:{33,33}]
  wire  _GEN_238 = 7'h6e == reqIndex ? way0V_110 : _GEN_237; // @[ICache.scala 48:{33,33}]
  wire  _GEN_239 = 7'h6f == reqIndex ? way0V_111 : _GEN_238; // @[ICache.scala 48:{33,33}]
  wire  _GEN_240 = 7'h70 == reqIndex ? way0V_112 : _GEN_239; // @[ICache.scala 48:{33,33}]
  wire  _GEN_241 = 7'h71 == reqIndex ? way0V_113 : _GEN_240; // @[ICache.scala 48:{33,33}]
  wire  _GEN_242 = 7'h72 == reqIndex ? way0V_114 : _GEN_241; // @[ICache.scala 48:{33,33}]
  wire  _GEN_243 = 7'h73 == reqIndex ? way0V_115 : _GEN_242; // @[ICache.scala 48:{33,33}]
  wire  _GEN_244 = 7'h74 == reqIndex ? way0V_116 : _GEN_243; // @[ICache.scala 48:{33,33}]
  wire  _GEN_245 = 7'h75 == reqIndex ? way0V_117 : _GEN_244; // @[ICache.scala 48:{33,33}]
  wire  _GEN_246 = 7'h76 == reqIndex ? way0V_118 : _GEN_245; // @[ICache.scala 48:{33,33}]
  wire  _GEN_247 = 7'h77 == reqIndex ? way0V_119 : _GEN_246; // @[ICache.scala 48:{33,33}]
  wire  _GEN_248 = 7'h78 == reqIndex ? way0V_120 : _GEN_247; // @[ICache.scala 48:{33,33}]
  wire  _GEN_249 = 7'h79 == reqIndex ? way0V_121 : _GEN_248; // @[ICache.scala 48:{33,33}]
  wire  _GEN_250 = 7'h7a == reqIndex ? way0V_122 : _GEN_249; // @[ICache.scala 48:{33,33}]
  wire  _GEN_251 = 7'h7b == reqIndex ? way0V_123 : _GEN_250; // @[ICache.scala 48:{33,33}]
  wire  _GEN_252 = 7'h7c == reqIndex ? way0V_124 : _GEN_251; // @[ICache.scala 48:{33,33}]
  wire  _GEN_253 = 7'h7d == reqIndex ? way0V_125 : _GEN_252; // @[ICache.scala 48:{33,33}]
  wire  _GEN_254 = 7'h7e == reqIndex ? way0V_126 : _GEN_253; // @[ICache.scala 48:{33,33}]
  wire  _GEN_255 = 7'h7f == reqIndex ? way0V_127 : _GEN_254; // @[ICache.scala 48:{33,33}]
  wire  way0Hit = _GEN_255 & _GEN_127 == reqTag; // @[ICache.scala 48:33]
  wire [20:0] _GEN_257 = 7'h1 == reqIndex ? way1Tag_1 : way1Tag_0; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_258 = 7'h2 == reqIndex ? way1Tag_2 : _GEN_257; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_259 = 7'h3 == reqIndex ? way1Tag_3 : _GEN_258; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_260 = 7'h4 == reqIndex ? way1Tag_4 : _GEN_259; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_261 = 7'h5 == reqIndex ? way1Tag_5 : _GEN_260; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_262 = 7'h6 == reqIndex ? way1Tag_6 : _GEN_261; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_263 = 7'h7 == reqIndex ? way1Tag_7 : _GEN_262; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_264 = 7'h8 == reqIndex ? way1Tag_8 : _GEN_263; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_265 = 7'h9 == reqIndex ? way1Tag_9 : _GEN_264; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_266 = 7'ha == reqIndex ? way1Tag_10 : _GEN_265; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_267 = 7'hb == reqIndex ? way1Tag_11 : _GEN_266; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_268 = 7'hc == reqIndex ? way1Tag_12 : _GEN_267; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_269 = 7'hd == reqIndex ? way1Tag_13 : _GEN_268; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_270 = 7'he == reqIndex ? way1Tag_14 : _GEN_269; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_271 = 7'hf == reqIndex ? way1Tag_15 : _GEN_270; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_272 = 7'h10 == reqIndex ? way1Tag_16 : _GEN_271; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_273 = 7'h11 == reqIndex ? way1Tag_17 : _GEN_272; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_274 = 7'h12 == reqIndex ? way1Tag_18 : _GEN_273; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_275 = 7'h13 == reqIndex ? way1Tag_19 : _GEN_274; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_276 = 7'h14 == reqIndex ? way1Tag_20 : _GEN_275; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_277 = 7'h15 == reqIndex ? way1Tag_21 : _GEN_276; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_278 = 7'h16 == reqIndex ? way1Tag_22 : _GEN_277; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_279 = 7'h17 == reqIndex ? way1Tag_23 : _GEN_278; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_280 = 7'h18 == reqIndex ? way1Tag_24 : _GEN_279; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_281 = 7'h19 == reqIndex ? way1Tag_25 : _GEN_280; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_282 = 7'h1a == reqIndex ? way1Tag_26 : _GEN_281; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_283 = 7'h1b == reqIndex ? way1Tag_27 : _GEN_282; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_284 = 7'h1c == reqIndex ? way1Tag_28 : _GEN_283; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_285 = 7'h1d == reqIndex ? way1Tag_29 : _GEN_284; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_286 = 7'h1e == reqIndex ? way1Tag_30 : _GEN_285; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_287 = 7'h1f == reqIndex ? way1Tag_31 : _GEN_286; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_288 = 7'h20 == reqIndex ? way1Tag_32 : _GEN_287; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_289 = 7'h21 == reqIndex ? way1Tag_33 : _GEN_288; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_290 = 7'h22 == reqIndex ? way1Tag_34 : _GEN_289; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_291 = 7'h23 == reqIndex ? way1Tag_35 : _GEN_290; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_292 = 7'h24 == reqIndex ? way1Tag_36 : _GEN_291; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_293 = 7'h25 == reqIndex ? way1Tag_37 : _GEN_292; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_294 = 7'h26 == reqIndex ? way1Tag_38 : _GEN_293; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_295 = 7'h27 == reqIndex ? way1Tag_39 : _GEN_294; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_296 = 7'h28 == reqIndex ? way1Tag_40 : _GEN_295; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_297 = 7'h29 == reqIndex ? way1Tag_41 : _GEN_296; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_298 = 7'h2a == reqIndex ? way1Tag_42 : _GEN_297; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_299 = 7'h2b == reqIndex ? way1Tag_43 : _GEN_298; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_300 = 7'h2c == reqIndex ? way1Tag_44 : _GEN_299; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_301 = 7'h2d == reqIndex ? way1Tag_45 : _GEN_300; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_302 = 7'h2e == reqIndex ? way1Tag_46 : _GEN_301; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_303 = 7'h2f == reqIndex ? way1Tag_47 : _GEN_302; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_304 = 7'h30 == reqIndex ? way1Tag_48 : _GEN_303; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_305 = 7'h31 == reqIndex ? way1Tag_49 : _GEN_304; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_306 = 7'h32 == reqIndex ? way1Tag_50 : _GEN_305; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_307 = 7'h33 == reqIndex ? way1Tag_51 : _GEN_306; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_308 = 7'h34 == reqIndex ? way1Tag_52 : _GEN_307; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_309 = 7'h35 == reqIndex ? way1Tag_53 : _GEN_308; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_310 = 7'h36 == reqIndex ? way1Tag_54 : _GEN_309; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_311 = 7'h37 == reqIndex ? way1Tag_55 : _GEN_310; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_312 = 7'h38 == reqIndex ? way1Tag_56 : _GEN_311; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_313 = 7'h39 == reqIndex ? way1Tag_57 : _GEN_312; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_314 = 7'h3a == reqIndex ? way1Tag_58 : _GEN_313; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_315 = 7'h3b == reqIndex ? way1Tag_59 : _GEN_314; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_316 = 7'h3c == reqIndex ? way1Tag_60 : _GEN_315; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_317 = 7'h3d == reqIndex ? way1Tag_61 : _GEN_316; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_318 = 7'h3e == reqIndex ? way1Tag_62 : _GEN_317; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_319 = 7'h3f == reqIndex ? way1Tag_63 : _GEN_318; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_320 = 7'h40 == reqIndex ? way1Tag_64 : _GEN_319; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_321 = 7'h41 == reqIndex ? way1Tag_65 : _GEN_320; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_322 = 7'h42 == reqIndex ? way1Tag_66 : _GEN_321; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_323 = 7'h43 == reqIndex ? way1Tag_67 : _GEN_322; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_324 = 7'h44 == reqIndex ? way1Tag_68 : _GEN_323; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_325 = 7'h45 == reqIndex ? way1Tag_69 : _GEN_324; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_326 = 7'h46 == reqIndex ? way1Tag_70 : _GEN_325; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_327 = 7'h47 == reqIndex ? way1Tag_71 : _GEN_326; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_328 = 7'h48 == reqIndex ? way1Tag_72 : _GEN_327; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_329 = 7'h49 == reqIndex ? way1Tag_73 : _GEN_328; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_330 = 7'h4a == reqIndex ? way1Tag_74 : _GEN_329; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_331 = 7'h4b == reqIndex ? way1Tag_75 : _GEN_330; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_332 = 7'h4c == reqIndex ? way1Tag_76 : _GEN_331; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_333 = 7'h4d == reqIndex ? way1Tag_77 : _GEN_332; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_334 = 7'h4e == reqIndex ? way1Tag_78 : _GEN_333; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_335 = 7'h4f == reqIndex ? way1Tag_79 : _GEN_334; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_336 = 7'h50 == reqIndex ? way1Tag_80 : _GEN_335; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_337 = 7'h51 == reqIndex ? way1Tag_81 : _GEN_336; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_338 = 7'h52 == reqIndex ? way1Tag_82 : _GEN_337; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_339 = 7'h53 == reqIndex ? way1Tag_83 : _GEN_338; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_340 = 7'h54 == reqIndex ? way1Tag_84 : _GEN_339; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_341 = 7'h55 == reqIndex ? way1Tag_85 : _GEN_340; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_342 = 7'h56 == reqIndex ? way1Tag_86 : _GEN_341; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_343 = 7'h57 == reqIndex ? way1Tag_87 : _GEN_342; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_344 = 7'h58 == reqIndex ? way1Tag_88 : _GEN_343; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_345 = 7'h59 == reqIndex ? way1Tag_89 : _GEN_344; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_346 = 7'h5a == reqIndex ? way1Tag_90 : _GEN_345; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_347 = 7'h5b == reqIndex ? way1Tag_91 : _GEN_346; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_348 = 7'h5c == reqIndex ? way1Tag_92 : _GEN_347; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_349 = 7'h5d == reqIndex ? way1Tag_93 : _GEN_348; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_350 = 7'h5e == reqIndex ? way1Tag_94 : _GEN_349; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_351 = 7'h5f == reqIndex ? way1Tag_95 : _GEN_350; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_352 = 7'h60 == reqIndex ? way1Tag_96 : _GEN_351; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_353 = 7'h61 == reqIndex ? way1Tag_97 : _GEN_352; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_354 = 7'h62 == reqIndex ? way1Tag_98 : _GEN_353; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_355 = 7'h63 == reqIndex ? way1Tag_99 : _GEN_354; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_356 = 7'h64 == reqIndex ? way1Tag_100 : _GEN_355; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_357 = 7'h65 == reqIndex ? way1Tag_101 : _GEN_356; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_358 = 7'h66 == reqIndex ? way1Tag_102 : _GEN_357; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_359 = 7'h67 == reqIndex ? way1Tag_103 : _GEN_358; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_360 = 7'h68 == reqIndex ? way1Tag_104 : _GEN_359; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_361 = 7'h69 == reqIndex ? way1Tag_105 : _GEN_360; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_362 = 7'h6a == reqIndex ? way1Tag_106 : _GEN_361; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_363 = 7'h6b == reqIndex ? way1Tag_107 : _GEN_362; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_364 = 7'h6c == reqIndex ? way1Tag_108 : _GEN_363; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_365 = 7'h6d == reqIndex ? way1Tag_109 : _GEN_364; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_366 = 7'h6e == reqIndex ? way1Tag_110 : _GEN_365; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_367 = 7'h6f == reqIndex ? way1Tag_111 : _GEN_366; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_368 = 7'h70 == reqIndex ? way1Tag_112 : _GEN_367; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_369 = 7'h71 == reqIndex ? way1Tag_113 : _GEN_368; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_370 = 7'h72 == reqIndex ? way1Tag_114 : _GEN_369; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_371 = 7'h73 == reqIndex ? way1Tag_115 : _GEN_370; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_372 = 7'h74 == reqIndex ? way1Tag_116 : _GEN_371; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_373 = 7'h75 == reqIndex ? way1Tag_117 : _GEN_372; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_374 = 7'h76 == reqIndex ? way1Tag_118 : _GEN_373; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_375 = 7'h77 == reqIndex ? way1Tag_119 : _GEN_374; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_376 = 7'h78 == reqIndex ? way1Tag_120 : _GEN_375; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_377 = 7'h79 == reqIndex ? way1Tag_121 : _GEN_376; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_378 = 7'h7a == reqIndex ? way1Tag_122 : _GEN_377; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_379 = 7'h7b == reqIndex ? way1Tag_123 : _GEN_378; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_380 = 7'h7c == reqIndex ? way1Tag_124 : _GEN_379; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_381 = 7'h7d == reqIndex ? way1Tag_125 : _GEN_380; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_382 = 7'h7e == reqIndex ? way1Tag_126 : _GEN_381; // @[ICache.scala 49:{55,55}]
  wire [20:0] _GEN_383 = 7'h7f == reqIndex ? way1Tag_127 : _GEN_382; // @[ICache.scala 49:{55,55}]
  wire  _GEN_385 = 7'h1 == reqIndex ? way1V_1 : way1V_0; // @[ICache.scala 49:{33,33}]
  wire  _GEN_386 = 7'h2 == reqIndex ? way1V_2 : _GEN_385; // @[ICache.scala 49:{33,33}]
  wire  _GEN_387 = 7'h3 == reqIndex ? way1V_3 : _GEN_386; // @[ICache.scala 49:{33,33}]
  wire  _GEN_388 = 7'h4 == reqIndex ? way1V_4 : _GEN_387; // @[ICache.scala 49:{33,33}]
  wire  _GEN_389 = 7'h5 == reqIndex ? way1V_5 : _GEN_388; // @[ICache.scala 49:{33,33}]
  wire  _GEN_390 = 7'h6 == reqIndex ? way1V_6 : _GEN_389; // @[ICache.scala 49:{33,33}]
  wire  _GEN_391 = 7'h7 == reqIndex ? way1V_7 : _GEN_390; // @[ICache.scala 49:{33,33}]
  wire  _GEN_392 = 7'h8 == reqIndex ? way1V_8 : _GEN_391; // @[ICache.scala 49:{33,33}]
  wire  _GEN_393 = 7'h9 == reqIndex ? way1V_9 : _GEN_392; // @[ICache.scala 49:{33,33}]
  wire  _GEN_394 = 7'ha == reqIndex ? way1V_10 : _GEN_393; // @[ICache.scala 49:{33,33}]
  wire  _GEN_395 = 7'hb == reqIndex ? way1V_11 : _GEN_394; // @[ICache.scala 49:{33,33}]
  wire  _GEN_396 = 7'hc == reqIndex ? way1V_12 : _GEN_395; // @[ICache.scala 49:{33,33}]
  wire  _GEN_397 = 7'hd == reqIndex ? way1V_13 : _GEN_396; // @[ICache.scala 49:{33,33}]
  wire  _GEN_398 = 7'he == reqIndex ? way1V_14 : _GEN_397; // @[ICache.scala 49:{33,33}]
  wire  _GEN_399 = 7'hf == reqIndex ? way1V_15 : _GEN_398; // @[ICache.scala 49:{33,33}]
  wire  _GEN_400 = 7'h10 == reqIndex ? way1V_16 : _GEN_399; // @[ICache.scala 49:{33,33}]
  wire  _GEN_401 = 7'h11 == reqIndex ? way1V_17 : _GEN_400; // @[ICache.scala 49:{33,33}]
  wire  _GEN_402 = 7'h12 == reqIndex ? way1V_18 : _GEN_401; // @[ICache.scala 49:{33,33}]
  wire  _GEN_403 = 7'h13 == reqIndex ? way1V_19 : _GEN_402; // @[ICache.scala 49:{33,33}]
  wire  _GEN_404 = 7'h14 == reqIndex ? way1V_20 : _GEN_403; // @[ICache.scala 49:{33,33}]
  wire  _GEN_405 = 7'h15 == reqIndex ? way1V_21 : _GEN_404; // @[ICache.scala 49:{33,33}]
  wire  _GEN_406 = 7'h16 == reqIndex ? way1V_22 : _GEN_405; // @[ICache.scala 49:{33,33}]
  wire  _GEN_407 = 7'h17 == reqIndex ? way1V_23 : _GEN_406; // @[ICache.scala 49:{33,33}]
  wire  _GEN_408 = 7'h18 == reqIndex ? way1V_24 : _GEN_407; // @[ICache.scala 49:{33,33}]
  wire  _GEN_409 = 7'h19 == reqIndex ? way1V_25 : _GEN_408; // @[ICache.scala 49:{33,33}]
  wire  _GEN_410 = 7'h1a == reqIndex ? way1V_26 : _GEN_409; // @[ICache.scala 49:{33,33}]
  wire  _GEN_411 = 7'h1b == reqIndex ? way1V_27 : _GEN_410; // @[ICache.scala 49:{33,33}]
  wire  _GEN_412 = 7'h1c == reqIndex ? way1V_28 : _GEN_411; // @[ICache.scala 49:{33,33}]
  wire  _GEN_413 = 7'h1d == reqIndex ? way1V_29 : _GEN_412; // @[ICache.scala 49:{33,33}]
  wire  _GEN_414 = 7'h1e == reqIndex ? way1V_30 : _GEN_413; // @[ICache.scala 49:{33,33}]
  wire  _GEN_415 = 7'h1f == reqIndex ? way1V_31 : _GEN_414; // @[ICache.scala 49:{33,33}]
  wire  _GEN_416 = 7'h20 == reqIndex ? way1V_32 : _GEN_415; // @[ICache.scala 49:{33,33}]
  wire  _GEN_417 = 7'h21 == reqIndex ? way1V_33 : _GEN_416; // @[ICache.scala 49:{33,33}]
  wire  _GEN_418 = 7'h22 == reqIndex ? way1V_34 : _GEN_417; // @[ICache.scala 49:{33,33}]
  wire  _GEN_419 = 7'h23 == reqIndex ? way1V_35 : _GEN_418; // @[ICache.scala 49:{33,33}]
  wire  _GEN_420 = 7'h24 == reqIndex ? way1V_36 : _GEN_419; // @[ICache.scala 49:{33,33}]
  wire  _GEN_421 = 7'h25 == reqIndex ? way1V_37 : _GEN_420; // @[ICache.scala 49:{33,33}]
  wire  _GEN_422 = 7'h26 == reqIndex ? way1V_38 : _GEN_421; // @[ICache.scala 49:{33,33}]
  wire  _GEN_423 = 7'h27 == reqIndex ? way1V_39 : _GEN_422; // @[ICache.scala 49:{33,33}]
  wire  _GEN_424 = 7'h28 == reqIndex ? way1V_40 : _GEN_423; // @[ICache.scala 49:{33,33}]
  wire  _GEN_425 = 7'h29 == reqIndex ? way1V_41 : _GEN_424; // @[ICache.scala 49:{33,33}]
  wire  _GEN_426 = 7'h2a == reqIndex ? way1V_42 : _GEN_425; // @[ICache.scala 49:{33,33}]
  wire  _GEN_427 = 7'h2b == reqIndex ? way1V_43 : _GEN_426; // @[ICache.scala 49:{33,33}]
  wire  _GEN_428 = 7'h2c == reqIndex ? way1V_44 : _GEN_427; // @[ICache.scala 49:{33,33}]
  wire  _GEN_429 = 7'h2d == reqIndex ? way1V_45 : _GEN_428; // @[ICache.scala 49:{33,33}]
  wire  _GEN_430 = 7'h2e == reqIndex ? way1V_46 : _GEN_429; // @[ICache.scala 49:{33,33}]
  wire  _GEN_431 = 7'h2f == reqIndex ? way1V_47 : _GEN_430; // @[ICache.scala 49:{33,33}]
  wire  _GEN_432 = 7'h30 == reqIndex ? way1V_48 : _GEN_431; // @[ICache.scala 49:{33,33}]
  wire  _GEN_433 = 7'h31 == reqIndex ? way1V_49 : _GEN_432; // @[ICache.scala 49:{33,33}]
  wire  _GEN_434 = 7'h32 == reqIndex ? way1V_50 : _GEN_433; // @[ICache.scala 49:{33,33}]
  wire  _GEN_435 = 7'h33 == reqIndex ? way1V_51 : _GEN_434; // @[ICache.scala 49:{33,33}]
  wire  _GEN_436 = 7'h34 == reqIndex ? way1V_52 : _GEN_435; // @[ICache.scala 49:{33,33}]
  wire  _GEN_437 = 7'h35 == reqIndex ? way1V_53 : _GEN_436; // @[ICache.scala 49:{33,33}]
  wire  _GEN_438 = 7'h36 == reqIndex ? way1V_54 : _GEN_437; // @[ICache.scala 49:{33,33}]
  wire  _GEN_439 = 7'h37 == reqIndex ? way1V_55 : _GEN_438; // @[ICache.scala 49:{33,33}]
  wire  _GEN_440 = 7'h38 == reqIndex ? way1V_56 : _GEN_439; // @[ICache.scala 49:{33,33}]
  wire  _GEN_441 = 7'h39 == reqIndex ? way1V_57 : _GEN_440; // @[ICache.scala 49:{33,33}]
  wire  _GEN_442 = 7'h3a == reqIndex ? way1V_58 : _GEN_441; // @[ICache.scala 49:{33,33}]
  wire  _GEN_443 = 7'h3b == reqIndex ? way1V_59 : _GEN_442; // @[ICache.scala 49:{33,33}]
  wire  _GEN_444 = 7'h3c == reqIndex ? way1V_60 : _GEN_443; // @[ICache.scala 49:{33,33}]
  wire  _GEN_445 = 7'h3d == reqIndex ? way1V_61 : _GEN_444; // @[ICache.scala 49:{33,33}]
  wire  _GEN_446 = 7'h3e == reqIndex ? way1V_62 : _GEN_445; // @[ICache.scala 49:{33,33}]
  wire  _GEN_447 = 7'h3f == reqIndex ? way1V_63 : _GEN_446; // @[ICache.scala 49:{33,33}]
  wire  _GEN_448 = 7'h40 == reqIndex ? way1V_64 : _GEN_447; // @[ICache.scala 49:{33,33}]
  wire  _GEN_449 = 7'h41 == reqIndex ? way1V_65 : _GEN_448; // @[ICache.scala 49:{33,33}]
  wire  _GEN_450 = 7'h42 == reqIndex ? way1V_66 : _GEN_449; // @[ICache.scala 49:{33,33}]
  wire  _GEN_451 = 7'h43 == reqIndex ? way1V_67 : _GEN_450; // @[ICache.scala 49:{33,33}]
  wire  _GEN_452 = 7'h44 == reqIndex ? way1V_68 : _GEN_451; // @[ICache.scala 49:{33,33}]
  wire  _GEN_453 = 7'h45 == reqIndex ? way1V_69 : _GEN_452; // @[ICache.scala 49:{33,33}]
  wire  _GEN_454 = 7'h46 == reqIndex ? way1V_70 : _GEN_453; // @[ICache.scala 49:{33,33}]
  wire  _GEN_455 = 7'h47 == reqIndex ? way1V_71 : _GEN_454; // @[ICache.scala 49:{33,33}]
  wire  _GEN_456 = 7'h48 == reqIndex ? way1V_72 : _GEN_455; // @[ICache.scala 49:{33,33}]
  wire  _GEN_457 = 7'h49 == reqIndex ? way1V_73 : _GEN_456; // @[ICache.scala 49:{33,33}]
  wire  _GEN_458 = 7'h4a == reqIndex ? way1V_74 : _GEN_457; // @[ICache.scala 49:{33,33}]
  wire  _GEN_459 = 7'h4b == reqIndex ? way1V_75 : _GEN_458; // @[ICache.scala 49:{33,33}]
  wire  _GEN_460 = 7'h4c == reqIndex ? way1V_76 : _GEN_459; // @[ICache.scala 49:{33,33}]
  wire  _GEN_461 = 7'h4d == reqIndex ? way1V_77 : _GEN_460; // @[ICache.scala 49:{33,33}]
  wire  _GEN_462 = 7'h4e == reqIndex ? way1V_78 : _GEN_461; // @[ICache.scala 49:{33,33}]
  wire  _GEN_463 = 7'h4f == reqIndex ? way1V_79 : _GEN_462; // @[ICache.scala 49:{33,33}]
  wire  _GEN_464 = 7'h50 == reqIndex ? way1V_80 : _GEN_463; // @[ICache.scala 49:{33,33}]
  wire  _GEN_465 = 7'h51 == reqIndex ? way1V_81 : _GEN_464; // @[ICache.scala 49:{33,33}]
  wire  _GEN_466 = 7'h52 == reqIndex ? way1V_82 : _GEN_465; // @[ICache.scala 49:{33,33}]
  wire  _GEN_467 = 7'h53 == reqIndex ? way1V_83 : _GEN_466; // @[ICache.scala 49:{33,33}]
  wire  _GEN_468 = 7'h54 == reqIndex ? way1V_84 : _GEN_467; // @[ICache.scala 49:{33,33}]
  wire  _GEN_469 = 7'h55 == reqIndex ? way1V_85 : _GEN_468; // @[ICache.scala 49:{33,33}]
  wire  _GEN_470 = 7'h56 == reqIndex ? way1V_86 : _GEN_469; // @[ICache.scala 49:{33,33}]
  wire  _GEN_471 = 7'h57 == reqIndex ? way1V_87 : _GEN_470; // @[ICache.scala 49:{33,33}]
  wire  _GEN_472 = 7'h58 == reqIndex ? way1V_88 : _GEN_471; // @[ICache.scala 49:{33,33}]
  wire  _GEN_473 = 7'h59 == reqIndex ? way1V_89 : _GEN_472; // @[ICache.scala 49:{33,33}]
  wire  _GEN_474 = 7'h5a == reqIndex ? way1V_90 : _GEN_473; // @[ICache.scala 49:{33,33}]
  wire  _GEN_475 = 7'h5b == reqIndex ? way1V_91 : _GEN_474; // @[ICache.scala 49:{33,33}]
  wire  _GEN_476 = 7'h5c == reqIndex ? way1V_92 : _GEN_475; // @[ICache.scala 49:{33,33}]
  wire  _GEN_477 = 7'h5d == reqIndex ? way1V_93 : _GEN_476; // @[ICache.scala 49:{33,33}]
  wire  _GEN_478 = 7'h5e == reqIndex ? way1V_94 : _GEN_477; // @[ICache.scala 49:{33,33}]
  wire  _GEN_479 = 7'h5f == reqIndex ? way1V_95 : _GEN_478; // @[ICache.scala 49:{33,33}]
  wire  _GEN_480 = 7'h60 == reqIndex ? way1V_96 : _GEN_479; // @[ICache.scala 49:{33,33}]
  wire  _GEN_481 = 7'h61 == reqIndex ? way1V_97 : _GEN_480; // @[ICache.scala 49:{33,33}]
  wire  _GEN_482 = 7'h62 == reqIndex ? way1V_98 : _GEN_481; // @[ICache.scala 49:{33,33}]
  wire  _GEN_483 = 7'h63 == reqIndex ? way1V_99 : _GEN_482; // @[ICache.scala 49:{33,33}]
  wire  _GEN_484 = 7'h64 == reqIndex ? way1V_100 : _GEN_483; // @[ICache.scala 49:{33,33}]
  wire  _GEN_485 = 7'h65 == reqIndex ? way1V_101 : _GEN_484; // @[ICache.scala 49:{33,33}]
  wire  _GEN_486 = 7'h66 == reqIndex ? way1V_102 : _GEN_485; // @[ICache.scala 49:{33,33}]
  wire  _GEN_487 = 7'h67 == reqIndex ? way1V_103 : _GEN_486; // @[ICache.scala 49:{33,33}]
  wire  _GEN_488 = 7'h68 == reqIndex ? way1V_104 : _GEN_487; // @[ICache.scala 49:{33,33}]
  wire  _GEN_489 = 7'h69 == reqIndex ? way1V_105 : _GEN_488; // @[ICache.scala 49:{33,33}]
  wire  _GEN_490 = 7'h6a == reqIndex ? way1V_106 : _GEN_489; // @[ICache.scala 49:{33,33}]
  wire  _GEN_491 = 7'h6b == reqIndex ? way1V_107 : _GEN_490; // @[ICache.scala 49:{33,33}]
  wire  _GEN_492 = 7'h6c == reqIndex ? way1V_108 : _GEN_491; // @[ICache.scala 49:{33,33}]
  wire  _GEN_493 = 7'h6d == reqIndex ? way1V_109 : _GEN_492; // @[ICache.scala 49:{33,33}]
  wire  _GEN_494 = 7'h6e == reqIndex ? way1V_110 : _GEN_493; // @[ICache.scala 49:{33,33}]
  wire  _GEN_495 = 7'h6f == reqIndex ? way1V_111 : _GEN_494; // @[ICache.scala 49:{33,33}]
  wire  _GEN_496 = 7'h70 == reqIndex ? way1V_112 : _GEN_495; // @[ICache.scala 49:{33,33}]
  wire  _GEN_497 = 7'h71 == reqIndex ? way1V_113 : _GEN_496; // @[ICache.scala 49:{33,33}]
  wire  _GEN_498 = 7'h72 == reqIndex ? way1V_114 : _GEN_497; // @[ICache.scala 49:{33,33}]
  wire  _GEN_499 = 7'h73 == reqIndex ? way1V_115 : _GEN_498; // @[ICache.scala 49:{33,33}]
  wire  _GEN_500 = 7'h74 == reqIndex ? way1V_116 : _GEN_499; // @[ICache.scala 49:{33,33}]
  wire  _GEN_501 = 7'h75 == reqIndex ? way1V_117 : _GEN_500; // @[ICache.scala 49:{33,33}]
  wire  _GEN_502 = 7'h76 == reqIndex ? way1V_118 : _GEN_501; // @[ICache.scala 49:{33,33}]
  wire  _GEN_503 = 7'h77 == reqIndex ? way1V_119 : _GEN_502; // @[ICache.scala 49:{33,33}]
  wire  _GEN_504 = 7'h78 == reqIndex ? way1V_120 : _GEN_503; // @[ICache.scala 49:{33,33}]
  wire  _GEN_505 = 7'h79 == reqIndex ? way1V_121 : _GEN_504; // @[ICache.scala 49:{33,33}]
  wire  _GEN_506 = 7'h7a == reqIndex ? way1V_122 : _GEN_505; // @[ICache.scala 49:{33,33}]
  wire  _GEN_507 = 7'h7b == reqIndex ? way1V_123 : _GEN_506; // @[ICache.scala 49:{33,33}]
  wire  _GEN_508 = 7'h7c == reqIndex ? way1V_124 : _GEN_507; // @[ICache.scala 49:{33,33}]
  wire  _GEN_509 = 7'h7d == reqIndex ? way1V_125 : _GEN_508; // @[ICache.scala 49:{33,33}]
  wire  _GEN_510 = 7'h7e == reqIndex ? way1V_126 : _GEN_509; // @[ICache.scala 49:{33,33}]
  wire  _GEN_511 = 7'h7f == reqIndex ? way1V_127 : _GEN_510; // @[ICache.scala 49:{33,33}]
  wire  way1Hit = _GEN_511 & _GEN_383 == reqTag; // @[ICache.scala 49:33]
  wire [7:0] _cacheRIndex_T = {1'h0,reqIndex}; // @[Cat.scala 31:58]
  wire [7:0] _cacheRIndex_T_1 = {1'h1,reqIndex}; // @[Cat.scala 31:58]
  wire [7:0] cacheRIndex = way0Hit ? _cacheRIndex_T : _cacheRIndex_T_1; // @[ICache.scala 50:24]
  wire  cacheHitEn = way0Hit | way1Hit; // @[ICache.scala 52:28]
  wire  sFillEn = state == 2'h3; // @[ICache.scala 108:23]
  wire  _GEN_520 = 7'h1 == reqIndex ? way0Age_1 : way0Age_0; // @[ICache.scala 110:{38,38}]
  wire  _GEN_521 = 7'h2 == reqIndex ? way0Age_2 : _GEN_520; // @[ICache.scala 110:{38,38}]
  wire  _GEN_522 = 7'h3 == reqIndex ? way0Age_3 : _GEN_521; // @[ICache.scala 110:{38,38}]
  wire  _GEN_523 = 7'h4 == reqIndex ? way0Age_4 : _GEN_522; // @[ICache.scala 110:{38,38}]
  wire  _GEN_524 = 7'h5 == reqIndex ? way0Age_5 : _GEN_523; // @[ICache.scala 110:{38,38}]
  wire  _GEN_525 = 7'h6 == reqIndex ? way0Age_6 : _GEN_524; // @[ICache.scala 110:{38,38}]
  wire  _GEN_526 = 7'h7 == reqIndex ? way0Age_7 : _GEN_525; // @[ICache.scala 110:{38,38}]
  wire  _GEN_527 = 7'h8 == reqIndex ? way0Age_8 : _GEN_526; // @[ICache.scala 110:{38,38}]
  wire  _GEN_528 = 7'h9 == reqIndex ? way0Age_9 : _GEN_527; // @[ICache.scala 110:{38,38}]
  wire  _GEN_529 = 7'ha == reqIndex ? way0Age_10 : _GEN_528; // @[ICache.scala 110:{38,38}]
  wire  _GEN_530 = 7'hb == reqIndex ? way0Age_11 : _GEN_529; // @[ICache.scala 110:{38,38}]
  wire  _GEN_531 = 7'hc == reqIndex ? way0Age_12 : _GEN_530; // @[ICache.scala 110:{38,38}]
  wire  _GEN_532 = 7'hd == reqIndex ? way0Age_13 : _GEN_531; // @[ICache.scala 110:{38,38}]
  wire  _GEN_533 = 7'he == reqIndex ? way0Age_14 : _GEN_532; // @[ICache.scala 110:{38,38}]
  wire  _GEN_534 = 7'hf == reqIndex ? way0Age_15 : _GEN_533; // @[ICache.scala 110:{38,38}]
  wire  _GEN_535 = 7'h10 == reqIndex ? way0Age_16 : _GEN_534; // @[ICache.scala 110:{38,38}]
  wire  _GEN_536 = 7'h11 == reqIndex ? way0Age_17 : _GEN_535; // @[ICache.scala 110:{38,38}]
  wire  _GEN_537 = 7'h12 == reqIndex ? way0Age_18 : _GEN_536; // @[ICache.scala 110:{38,38}]
  wire  _GEN_538 = 7'h13 == reqIndex ? way0Age_19 : _GEN_537; // @[ICache.scala 110:{38,38}]
  wire  _GEN_539 = 7'h14 == reqIndex ? way0Age_20 : _GEN_538; // @[ICache.scala 110:{38,38}]
  wire  _GEN_540 = 7'h15 == reqIndex ? way0Age_21 : _GEN_539; // @[ICache.scala 110:{38,38}]
  wire  _GEN_541 = 7'h16 == reqIndex ? way0Age_22 : _GEN_540; // @[ICache.scala 110:{38,38}]
  wire  _GEN_542 = 7'h17 == reqIndex ? way0Age_23 : _GEN_541; // @[ICache.scala 110:{38,38}]
  wire  _GEN_543 = 7'h18 == reqIndex ? way0Age_24 : _GEN_542; // @[ICache.scala 110:{38,38}]
  wire  _GEN_544 = 7'h19 == reqIndex ? way0Age_25 : _GEN_543; // @[ICache.scala 110:{38,38}]
  wire  _GEN_545 = 7'h1a == reqIndex ? way0Age_26 : _GEN_544; // @[ICache.scala 110:{38,38}]
  wire  _GEN_546 = 7'h1b == reqIndex ? way0Age_27 : _GEN_545; // @[ICache.scala 110:{38,38}]
  wire  _GEN_547 = 7'h1c == reqIndex ? way0Age_28 : _GEN_546; // @[ICache.scala 110:{38,38}]
  wire  _GEN_548 = 7'h1d == reqIndex ? way0Age_29 : _GEN_547; // @[ICache.scala 110:{38,38}]
  wire  _GEN_549 = 7'h1e == reqIndex ? way0Age_30 : _GEN_548; // @[ICache.scala 110:{38,38}]
  wire  _GEN_550 = 7'h1f == reqIndex ? way0Age_31 : _GEN_549; // @[ICache.scala 110:{38,38}]
  wire  _GEN_551 = 7'h20 == reqIndex ? way0Age_32 : _GEN_550; // @[ICache.scala 110:{38,38}]
  wire  _GEN_552 = 7'h21 == reqIndex ? way0Age_33 : _GEN_551; // @[ICache.scala 110:{38,38}]
  wire  _GEN_553 = 7'h22 == reqIndex ? way0Age_34 : _GEN_552; // @[ICache.scala 110:{38,38}]
  wire  _GEN_554 = 7'h23 == reqIndex ? way0Age_35 : _GEN_553; // @[ICache.scala 110:{38,38}]
  wire  _GEN_555 = 7'h24 == reqIndex ? way0Age_36 : _GEN_554; // @[ICache.scala 110:{38,38}]
  wire  _GEN_556 = 7'h25 == reqIndex ? way0Age_37 : _GEN_555; // @[ICache.scala 110:{38,38}]
  wire  _GEN_557 = 7'h26 == reqIndex ? way0Age_38 : _GEN_556; // @[ICache.scala 110:{38,38}]
  wire  _GEN_558 = 7'h27 == reqIndex ? way0Age_39 : _GEN_557; // @[ICache.scala 110:{38,38}]
  wire  _GEN_559 = 7'h28 == reqIndex ? way0Age_40 : _GEN_558; // @[ICache.scala 110:{38,38}]
  wire  _GEN_560 = 7'h29 == reqIndex ? way0Age_41 : _GEN_559; // @[ICache.scala 110:{38,38}]
  wire  _GEN_561 = 7'h2a == reqIndex ? way0Age_42 : _GEN_560; // @[ICache.scala 110:{38,38}]
  wire  _GEN_562 = 7'h2b == reqIndex ? way0Age_43 : _GEN_561; // @[ICache.scala 110:{38,38}]
  wire  _GEN_563 = 7'h2c == reqIndex ? way0Age_44 : _GEN_562; // @[ICache.scala 110:{38,38}]
  wire  _GEN_564 = 7'h2d == reqIndex ? way0Age_45 : _GEN_563; // @[ICache.scala 110:{38,38}]
  wire  _GEN_565 = 7'h2e == reqIndex ? way0Age_46 : _GEN_564; // @[ICache.scala 110:{38,38}]
  wire  _GEN_566 = 7'h2f == reqIndex ? way0Age_47 : _GEN_565; // @[ICache.scala 110:{38,38}]
  wire  _GEN_567 = 7'h30 == reqIndex ? way0Age_48 : _GEN_566; // @[ICache.scala 110:{38,38}]
  wire  _GEN_568 = 7'h31 == reqIndex ? way0Age_49 : _GEN_567; // @[ICache.scala 110:{38,38}]
  wire  _GEN_569 = 7'h32 == reqIndex ? way0Age_50 : _GEN_568; // @[ICache.scala 110:{38,38}]
  wire  _GEN_570 = 7'h33 == reqIndex ? way0Age_51 : _GEN_569; // @[ICache.scala 110:{38,38}]
  wire  _GEN_571 = 7'h34 == reqIndex ? way0Age_52 : _GEN_570; // @[ICache.scala 110:{38,38}]
  wire  _GEN_572 = 7'h35 == reqIndex ? way0Age_53 : _GEN_571; // @[ICache.scala 110:{38,38}]
  wire  _GEN_573 = 7'h36 == reqIndex ? way0Age_54 : _GEN_572; // @[ICache.scala 110:{38,38}]
  wire  _GEN_574 = 7'h37 == reqIndex ? way0Age_55 : _GEN_573; // @[ICache.scala 110:{38,38}]
  wire  _GEN_575 = 7'h38 == reqIndex ? way0Age_56 : _GEN_574; // @[ICache.scala 110:{38,38}]
  wire  _GEN_576 = 7'h39 == reqIndex ? way0Age_57 : _GEN_575; // @[ICache.scala 110:{38,38}]
  wire  _GEN_577 = 7'h3a == reqIndex ? way0Age_58 : _GEN_576; // @[ICache.scala 110:{38,38}]
  wire  _GEN_578 = 7'h3b == reqIndex ? way0Age_59 : _GEN_577; // @[ICache.scala 110:{38,38}]
  wire  _GEN_579 = 7'h3c == reqIndex ? way0Age_60 : _GEN_578; // @[ICache.scala 110:{38,38}]
  wire  _GEN_580 = 7'h3d == reqIndex ? way0Age_61 : _GEN_579; // @[ICache.scala 110:{38,38}]
  wire  _GEN_581 = 7'h3e == reqIndex ? way0Age_62 : _GEN_580; // @[ICache.scala 110:{38,38}]
  wire  _GEN_582 = 7'h3f == reqIndex ? way0Age_63 : _GEN_581; // @[ICache.scala 110:{38,38}]
  wire  _GEN_583 = 7'h40 == reqIndex ? way0Age_64 : _GEN_582; // @[ICache.scala 110:{38,38}]
  wire  _GEN_584 = 7'h41 == reqIndex ? way0Age_65 : _GEN_583; // @[ICache.scala 110:{38,38}]
  wire  _GEN_585 = 7'h42 == reqIndex ? way0Age_66 : _GEN_584; // @[ICache.scala 110:{38,38}]
  wire  _GEN_586 = 7'h43 == reqIndex ? way0Age_67 : _GEN_585; // @[ICache.scala 110:{38,38}]
  wire  _GEN_587 = 7'h44 == reqIndex ? way0Age_68 : _GEN_586; // @[ICache.scala 110:{38,38}]
  wire  _GEN_588 = 7'h45 == reqIndex ? way0Age_69 : _GEN_587; // @[ICache.scala 110:{38,38}]
  wire  _GEN_589 = 7'h46 == reqIndex ? way0Age_70 : _GEN_588; // @[ICache.scala 110:{38,38}]
  wire  _GEN_590 = 7'h47 == reqIndex ? way0Age_71 : _GEN_589; // @[ICache.scala 110:{38,38}]
  wire  _GEN_591 = 7'h48 == reqIndex ? way0Age_72 : _GEN_590; // @[ICache.scala 110:{38,38}]
  wire  _GEN_592 = 7'h49 == reqIndex ? way0Age_73 : _GEN_591; // @[ICache.scala 110:{38,38}]
  wire  _GEN_593 = 7'h4a == reqIndex ? way0Age_74 : _GEN_592; // @[ICache.scala 110:{38,38}]
  wire  _GEN_594 = 7'h4b == reqIndex ? way0Age_75 : _GEN_593; // @[ICache.scala 110:{38,38}]
  wire  _GEN_595 = 7'h4c == reqIndex ? way0Age_76 : _GEN_594; // @[ICache.scala 110:{38,38}]
  wire  _GEN_596 = 7'h4d == reqIndex ? way0Age_77 : _GEN_595; // @[ICache.scala 110:{38,38}]
  wire  _GEN_597 = 7'h4e == reqIndex ? way0Age_78 : _GEN_596; // @[ICache.scala 110:{38,38}]
  wire  _GEN_598 = 7'h4f == reqIndex ? way0Age_79 : _GEN_597; // @[ICache.scala 110:{38,38}]
  wire  _GEN_599 = 7'h50 == reqIndex ? way0Age_80 : _GEN_598; // @[ICache.scala 110:{38,38}]
  wire  _GEN_600 = 7'h51 == reqIndex ? way0Age_81 : _GEN_599; // @[ICache.scala 110:{38,38}]
  wire  _GEN_601 = 7'h52 == reqIndex ? way0Age_82 : _GEN_600; // @[ICache.scala 110:{38,38}]
  wire  _GEN_602 = 7'h53 == reqIndex ? way0Age_83 : _GEN_601; // @[ICache.scala 110:{38,38}]
  wire  _GEN_603 = 7'h54 == reqIndex ? way0Age_84 : _GEN_602; // @[ICache.scala 110:{38,38}]
  wire  _GEN_604 = 7'h55 == reqIndex ? way0Age_85 : _GEN_603; // @[ICache.scala 110:{38,38}]
  wire  _GEN_605 = 7'h56 == reqIndex ? way0Age_86 : _GEN_604; // @[ICache.scala 110:{38,38}]
  wire  _GEN_606 = 7'h57 == reqIndex ? way0Age_87 : _GEN_605; // @[ICache.scala 110:{38,38}]
  wire  _GEN_607 = 7'h58 == reqIndex ? way0Age_88 : _GEN_606; // @[ICache.scala 110:{38,38}]
  wire  _GEN_608 = 7'h59 == reqIndex ? way0Age_89 : _GEN_607; // @[ICache.scala 110:{38,38}]
  wire  _GEN_609 = 7'h5a == reqIndex ? way0Age_90 : _GEN_608; // @[ICache.scala 110:{38,38}]
  wire  _GEN_610 = 7'h5b == reqIndex ? way0Age_91 : _GEN_609; // @[ICache.scala 110:{38,38}]
  wire  _GEN_611 = 7'h5c == reqIndex ? way0Age_92 : _GEN_610; // @[ICache.scala 110:{38,38}]
  wire  _GEN_612 = 7'h5d == reqIndex ? way0Age_93 : _GEN_611; // @[ICache.scala 110:{38,38}]
  wire  _GEN_613 = 7'h5e == reqIndex ? way0Age_94 : _GEN_612; // @[ICache.scala 110:{38,38}]
  wire  _GEN_614 = 7'h5f == reqIndex ? way0Age_95 : _GEN_613; // @[ICache.scala 110:{38,38}]
  wire  _GEN_615 = 7'h60 == reqIndex ? way0Age_96 : _GEN_614; // @[ICache.scala 110:{38,38}]
  wire  _GEN_616 = 7'h61 == reqIndex ? way0Age_97 : _GEN_615; // @[ICache.scala 110:{38,38}]
  wire  _GEN_617 = 7'h62 == reqIndex ? way0Age_98 : _GEN_616; // @[ICache.scala 110:{38,38}]
  wire  _GEN_618 = 7'h63 == reqIndex ? way0Age_99 : _GEN_617; // @[ICache.scala 110:{38,38}]
  wire  _GEN_619 = 7'h64 == reqIndex ? way0Age_100 : _GEN_618; // @[ICache.scala 110:{38,38}]
  wire  _GEN_620 = 7'h65 == reqIndex ? way0Age_101 : _GEN_619; // @[ICache.scala 110:{38,38}]
  wire  _GEN_621 = 7'h66 == reqIndex ? way0Age_102 : _GEN_620; // @[ICache.scala 110:{38,38}]
  wire  _GEN_622 = 7'h67 == reqIndex ? way0Age_103 : _GEN_621; // @[ICache.scala 110:{38,38}]
  wire  _GEN_623 = 7'h68 == reqIndex ? way0Age_104 : _GEN_622; // @[ICache.scala 110:{38,38}]
  wire  _GEN_624 = 7'h69 == reqIndex ? way0Age_105 : _GEN_623; // @[ICache.scala 110:{38,38}]
  wire  _GEN_625 = 7'h6a == reqIndex ? way0Age_106 : _GEN_624; // @[ICache.scala 110:{38,38}]
  wire  _GEN_626 = 7'h6b == reqIndex ? way0Age_107 : _GEN_625; // @[ICache.scala 110:{38,38}]
  wire  _GEN_627 = 7'h6c == reqIndex ? way0Age_108 : _GEN_626; // @[ICache.scala 110:{38,38}]
  wire  _GEN_628 = 7'h6d == reqIndex ? way0Age_109 : _GEN_627; // @[ICache.scala 110:{38,38}]
  wire  _GEN_629 = 7'h6e == reqIndex ? way0Age_110 : _GEN_628; // @[ICache.scala 110:{38,38}]
  wire  _GEN_630 = 7'h6f == reqIndex ? way0Age_111 : _GEN_629; // @[ICache.scala 110:{38,38}]
  wire  _GEN_631 = 7'h70 == reqIndex ? way0Age_112 : _GEN_630; // @[ICache.scala 110:{38,38}]
  wire  _GEN_632 = 7'h71 == reqIndex ? way0Age_113 : _GEN_631; // @[ICache.scala 110:{38,38}]
  wire  _GEN_633 = 7'h72 == reqIndex ? way0Age_114 : _GEN_632; // @[ICache.scala 110:{38,38}]
  wire  _GEN_634 = 7'h73 == reqIndex ? way0Age_115 : _GEN_633; // @[ICache.scala 110:{38,38}]
  wire  _GEN_635 = 7'h74 == reqIndex ? way0Age_116 : _GEN_634; // @[ICache.scala 110:{38,38}]
  wire  _GEN_636 = 7'h75 == reqIndex ? way0Age_117 : _GEN_635; // @[ICache.scala 110:{38,38}]
  wire  _GEN_637 = 7'h76 == reqIndex ? way0Age_118 : _GEN_636; // @[ICache.scala 110:{38,38}]
  wire  _GEN_638 = 7'h77 == reqIndex ? way0Age_119 : _GEN_637; // @[ICache.scala 110:{38,38}]
  wire  _GEN_639 = 7'h78 == reqIndex ? way0Age_120 : _GEN_638; // @[ICache.scala 110:{38,38}]
  wire  _GEN_640 = 7'h79 == reqIndex ? way0Age_121 : _GEN_639; // @[ICache.scala 110:{38,38}]
  wire  _GEN_641 = 7'h7a == reqIndex ? way0Age_122 : _GEN_640; // @[ICache.scala 110:{38,38}]
  wire  _GEN_642 = 7'h7b == reqIndex ? way0Age_123 : _GEN_641; // @[ICache.scala 110:{38,38}]
  wire  _GEN_643 = 7'h7c == reqIndex ? way0Age_124 : _GEN_642; // @[ICache.scala 110:{38,38}]
  wire  _GEN_644 = 7'h7d == reqIndex ? way0Age_125 : _GEN_643; // @[ICache.scala 110:{38,38}]
  wire  _GEN_645 = 7'h7e == reqIndex ? way0Age_126 : _GEN_644; // @[ICache.scala 110:{38,38}]
  wire  _GEN_646 = 7'h7f == reqIndex ? way0Age_127 : _GEN_645; // @[ICache.scala 110:{38,38}]
  wire  ageWay0En = ~_GEN_646 & sFillEn; // @[ICache.scala 110:47]
  wire  cacheLineWay = ageWay0En ? 1'h0 : 1'h1; // @[ICache.scala 112:25]
  wire [7:0] cacheWIndex = {cacheLineWay,reqIndex}; // @[Cat.scala 31:58]
  wire [1:0] _GEN_514 = io_out_inst_ready ? 2'h3 : state; // @[ICache.scala 79:28 80:15 38:22]
  wire [1:0] _GEN_515 = 2'h3 == state ? 2'h1 : state; // @[ICache.scala 63:17 85:15 38:22]
  wire  sReadEn = state == 2'h1; // @[ICache.scala 89:23]
  wire [127:0] cacheRData = req_Q;
  wire [127:0] rData = sReadEn & cacheHitEn ? cacheRData : 128'h0; // @[ICache.scala 90:18]
  wire [31:0] _io_imem_inst_read_T_6 = 2'h1 == reqOff[3:2] ? rData[63:32] : rData[31:0]; // @[Mux.scala 81:58]
  wire [31:0] _io_imem_inst_read_T_8 = 2'h2 == reqOff[3:2] ? rData[95:64] : _io_imem_inst_read_T_6; // @[Mux.scala 81:58]
  wire  sAxiEn = state == 2'h2; // @[ICache.scala 100:22]
  wire  _GEN_648 = 7'h1 == reqIndex ? way1Age_1 : way1Age_0; // @[ICache.scala 111:{38,38}]
  wire  _GEN_649 = 7'h2 == reqIndex ? way1Age_2 : _GEN_648; // @[ICache.scala 111:{38,38}]
  wire  _GEN_650 = 7'h3 == reqIndex ? way1Age_3 : _GEN_649; // @[ICache.scala 111:{38,38}]
  wire  _GEN_651 = 7'h4 == reqIndex ? way1Age_4 : _GEN_650; // @[ICache.scala 111:{38,38}]
  wire  _GEN_652 = 7'h5 == reqIndex ? way1Age_5 : _GEN_651; // @[ICache.scala 111:{38,38}]
  wire  _GEN_653 = 7'h6 == reqIndex ? way1Age_6 : _GEN_652; // @[ICache.scala 111:{38,38}]
  wire  _GEN_654 = 7'h7 == reqIndex ? way1Age_7 : _GEN_653; // @[ICache.scala 111:{38,38}]
  wire  _GEN_655 = 7'h8 == reqIndex ? way1Age_8 : _GEN_654; // @[ICache.scala 111:{38,38}]
  wire  _GEN_656 = 7'h9 == reqIndex ? way1Age_9 : _GEN_655; // @[ICache.scala 111:{38,38}]
  wire  _GEN_657 = 7'ha == reqIndex ? way1Age_10 : _GEN_656; // @[ICache.scala 111:{38,38}]
  wire  _GEN_658 = 7'hb == reqIndex ? way1Age_11 : _GEN_657; // @[ICache.scala 111:{38,38}]
  wire  _GEN_659 = 7'hc == reqIndex ? way1Age_12 : _GEN_658; // @[ICache.scala 111:{38,38}]
  wire  _GEN_660 = 7'hd == reqIndex ? way1Age_13 : _GEN_659; // @[ICache.scala 111:{38,38}]
  wire  _GEN_661 = 7'he == reqIndex ? way1Age_14 : _GEN_660; // @[ICache.scala 111:{38,38}]
  wire  _GEN_662 = 7'hf == reqIndex ? way1Age_15 : _GEN_661; // @[ICache.scala 111:{38,38}]
  wire  _GEN_663 = 7'h10 == reqIndex ? way1Age_16 : _GEN_662; // @[ICache.scala 111:{38,38}]
  wire  _GEN_664 = 7'h11 == reqIndex ? way1Age_17 : _GEN_663; // @[ICache.scala 111:{38,38}]
  wire  _GEN_665 = 7'h12 == reqIndex ? way1Age_18 : _GEN_664; // @[ICache.scala 111:{38,38}]
  wire  _GEN_666 = 7'h13 == reqIndex ? way1Age_19 : _GEN_665; // @[ICache.scala 111:{38,38}]
  wire  _GEN_667 = 7'h14 == reqIndex ? way1Age_20 : _GEN_666; // @[ICache.scala 111:{38,38}]
  wire  _GEN_668 = 7'h15 == reqIndex ? way1Age_21 : _GEN_667; // @[ICache.scala 111:{38,38}]
  wire  _GEN_669 = 7'h16 == reqIndex ? way1Age_22 : _GEN_668; // @[ICache.scala 111:{38,38}]
  wire  _GEN_670 = 7'h17 == reqIndex ? way1Age_23 : _GEN_669; // @[ICache.scala 111:{38,38}]
  wire  _GEN_671 = 7'h18 == reqIndex ? way1Age_24 : _GEN_670; // @[ICache.scala 111:{38,38}]
  wire  _GEN_672 = 7'h19 == reqIndex ? way1Age_25 : _GEN_671; // @[ICache.scala 111:{38,38}]
  wire  _GEN_673 = 7'h1a == reqIndex ? way1Age_26 : _GEN_672; // @[ICache.scala 111:{38,38}]
  wire  _GEN_674 = 7'h1b == reqIndex ? way1Age_27 : _GEN_673; // @[ICache.scala 111:{38,38}]
  wire  _GEN_675 = 7'h1c == reqIndex ? way1Age_28 : _GEN_674; // @[ICache.scala 111:{38,38}]
  wire  _GEN_676 = 7'h1d == reqIndex ? way1Age_29 : _GEN_675; // @[ICache.scala 111:{38,38}]
  wire  _GEN_677 = 7'h1e == reqIndex ? way1Age_30 : _GEN_676; // @[ICache.scala 111:{38,38}]
  wire  _GEN_678 = 7'h1f == reqIndex ? way1Age_31 : _GEN_677; // @[ICache.scala 111:{38,38}]
  wire  _GEN_679 = 7'h20 == reqIndex ? way1Age_32 : _GEN_678; // @[ICache.scala 111:{38,38}]
  wire  _GEN_680 = 7'h21 == reqIndex ? way1Age_33 : _GEN_679; // @[ICache.scala 111:{38,38}]
  wire  _GEN_681 = 7'h22 == reqIndex ? way1Age_34 : _GEN_680; // @[ICache.scala 111:{38,38}]
  wire  _GEN_682 = 7'h23 == reqIndex ? way1Age_35 : _GEN_681; // @[ICache.scala 111:{38,38}]
  wire  _GEN_683 = 7'h24 == reqIndex ? way1Age_36 : _GEN_682; // @[ICache.scala 111:{38,38}]
  wire  _GEN_684 = 7'h25 == reqIndex ? way1Age_37 : _GEN_683; // @[ICache.scala 111:{38,38}]
  wire  _GEN_685 = 7'h26 == reqIndex ? way1Age_38 : _GEN_684; // @[ICache.scala 111:{38,38}]
  wire  _GEN_686 = 7'h27 == reqIndex ? way1Age_39 : _GEN_685; // @[ICache.scala 111:{38,38}]
  wire  _GEN_687 = 7'h28 == reqIndex ? way1Age_40 : _GEN_686; // @[ICache.scala 111:{38,38}]
  wire  _GEN_688 = 7'h29 == reqIndex ? way1Age_41 : _GEN_687; // @[ICache.scala 111:{38,38}]
  wire  _GEN_689 = 7'h2a == reqIndex ? way1Age_42 : _GEN_688; // @[ICache.scala 111:{38,38}]
  wire  _GEN_690 = 7'h2b == reqIndex ? way1Age_43 : _GEN_689; // @[ICache.scala 111:{38,38}]
  wire  _GEN_691 = 7'h2c == reqIndex ? way1Age_44 : _GEN_690; // @[ICache.scala 111:{38,38}]
  wire  _GEN_692 = 7'h2d == reqIndex ? way1Age_45 : _GEN_691; // @[ICache.scala 111:{38,38}]
  wire  _GEN_693 = 7'h2e == reqIndex ? way1Age_46 : _GEN_692; // @[ICache.scala 111:{38,38}]
  wire  _GEN_694 = 7'h2f == reqIndex ? way1Age_47 : _GEN_693; // @[ICache.scala 111:{38,38}]
  wire  _GEN_695 = 7'h30 == reqIndex ? way1Age_48 : _GEN_694; // @[ICache.scala 111:{38,38}]
  wire  _GEN_696 = 7'h31 == reqIndex ? way1Age_49 : _GEN_695; // @[ICache.scala 111:{38,38}]
  wire  _GEN_697 = 7'h32 == reqIndex ? way1Age_50 : _GEN_696; // @[ICache.scala 111:{38,38}]
  wire  _GEN_698 = 7'h33 == reqIndex ? way1Age_51 : _GEN_697; // @[ICache.scala 111:{38,38}]
  wire  _GEN_699 = 7'h34 == reqIndex ? way1Age_52 : _GEN_698; // @[ICache.scala 111:{38,38}]
  wire  _GEN_700 = 7'h35 == reqIndex ? way1Age_53 : _GEN_699; // @[ICache.scala 111:{38,38}]
  wire  _GEN_701 = 7'h36 == reqIndex ? way1Age_54 : _GEN_700; // @[ICache.scala 111:{38,38}]
  wire  _GEN_702 = 7'h37 == reqIndex ? way1Age_55 : _GEN_701; // @[ICache.scala 111:{38,38}]
  wire  _GEN_703 = 7'h38 == reqIndex ? way1Age_56 : _GEN_702; // @[ICache.scala 111:{38,38}]
  wire  _GEN_704 = 7'h39 == reqIndex ? way1Age_57 : _GEN_703; // @[ICache.scala 111:{38,38}]
  wire  _GEN_705 = 7'h3a == reqIndex ? way1Age_58 : _GEN_704; // @[ICache.scala 111:{38,38}]
  wire  _GEN_706 = 7'h3b == reqIndex ? way1Age_59 : _GEN_705; // @[ICache.scala 111:{38,38}]
  wire  _GEN_707 = 7'h3c == reqIndex ? way1Age_60 : _GEN_706; // @[ICache.scala 111:{38,38}]
  wire  _GEN_708 = 7'h3d == reqIndex ? way1Age_61 : _GEN_707; // @[ICache.scala 111:{38,38}]
  wire  _GEN_709 = 7'h3e == reqIndex ? way1Age_62 : _GEN_708; // @[ICache.scala 111:{38,38}]
  wire  _GEN_710 = 7'h3f == reqIndex ? way1Age_63 : _GEN_709; // @[ICache.scala 111:{38,38}]
  wire  _GEN_711 = 7'h40 == reqIndex ? way1Age_64 : _GEN_710; // @[ICache.scala 111:{38,38}]
  wire  _GEN_712 = 7'h41 == reqIndex ? way1Age_65 : _GEN_711; // @[ICache.scala 111:{38,38}]
  wire  _GEN_713 = 7'h42 == reqIndex ? way1Age_66 : _GEN_712; // @[ICache.scala 111:{38,38}]
  wire  _GEN_714 = 7'h43 == reqIndex ? way1Age_67 : _GEN_713; // @[ICache.scala 111:{38,38}]
  wire  _GEN_715 = 7'h44 == reqIndex ? way1Age_68 : _GEN_714; // @[ICache.scala 111:{38,38}]
  wire  _GEN_716 = 7'h45 == reqIndex ? way1Age_69 : _GEN_715; // @[ICache.scala 111:{38,38}]
  wire  _GEN_717 = 7'h46 == reqIndex ? way1Age_70 : _GEN_716; // @[ICache.scala 111:{38,38}]
  wire  _GEN_718 = 7'h47 == reqIndex ? way1Age_71 : _GEN_717; // @[ICache.scala 111:{38,38}]
  wire  _GEN_719 = 7'h48 == reqIndex ? way1Age_72 : _GEN_718; // @[ICache.scala 111:{38,38}]
  wire  _GEN_720 = 7'h49 == reqIndex ? way1Age_73 : _GEN_719; // @[ICache.scala 111:{38,38}]
  wire  _GEN_721 = 7'h4a == reqIndex ? way1Age_74 : _GEN_720; // @[ICache.scala 111:{38,38}]
  wire  _GEN_722 = 7'h4b == reqIndex ? way1Age_75 : _GEN_721; // @[ICache.scala 111:{38,38}]
  wire  _GEN_723 = 7'h4c == reqIndex ? way1Age_76 : _GEN_722; // @[ICache.scala 111:{38,38}]
  wire  _GEN_724 = 7'h4d == reqIndex ? way1Age_77 : _GEN_723; // @[ICache.scala 111:{38,38}]
  wire  _GEN_725 = 7'h4e == reqIndex ? way1Age_78 : _GEN_724; // @[ICache.scala 111:{38,38}]
  wire  _GEN_726 = 7'h4f == reqIndex ? way1Age_79 : _GEN_725; // @[ICache.scala 111:{38,38}]
  wire  _GEN_727 = 7'h50 == reqIndex ? way1Age_80 : _GEN_726; // @[ICache.scala 111:{38,38}]
  wire  _GEN_728 = 7'h51 == reqIndex ? way1Age_81 : _GEN_727; // @[ICache.scala 111:{38,38}]
  wire  _GEN_729 = 7'h52 == reqIndex ? way1Age_82 : _GEN_728; // @[ICache.scala 111:{38,38}]
  wire  _GEN_730 = 7'h53 == reqIndex ? way1Age_83 : _GEN_729; // @[ICache.scala 111:{38,38}]
  wire  _GEN_731 = 7'h54 == reqIndex ? way1Age_84 : _GEN_730; // @[ICache.scala 111:{38,38}]
  wire  _GEN_732 = 7'h55 == reqIndex ? way1Age_85 : _GEN_731; // @[ICache.scala 111:{38,38}]
  wire  _GEN_733 = 7'h56 == reqIndex ? way1Age_86 : _GEN_732; // @[ICache.scala 111:{38,38}]
  wire  _GEN_734 = 7'h57 == reqIndex ? way1Age_87 : _GEN_733; // @[ICache.scala 111:{38,38}]
  wire  _GEN_735 = 7'h58 == reqIndex ? way1Age_88 : _GEN_734; // @[ICache.scala 111:{38,38}]
  wire  _GEN_736 = 7'h59 == reqIndex ? way1Age_89 : _GEN_735; // @[ICache.scala 111:{38,38}]
  wire  _GEN_737 = 7'h5a == reqIndex ? way1Age_90 : _GEN_736; // @[ICache.scala 111:{38,38}]
  wire  _GEN_738 = 7'h5b == reqIndex ? way1Age_91 : _GEN_737; // @[ICache.scala 111:{38,38}]
  wire  _GEN_739 = 7'h5c == reqIndex ? way1Age_92 : _GEN_738; // @[ICache.scala 111:{38,38}]
  wire  _GEN_740 = 7'h5d == reqIndex ? way1Age_93 : _GEN_739; // @[ICache.scala 111:{38,38}]
  wire  _GEN_741 = 7'h5e == reqIndex ? way1Age_94 : _GEN_740; // @[ICache.scala 111:{38,38}]
  wire  _GEN_742 = 7'h5f == reqIndex ? way1Age_95 : _GEN_741; // @[ICache.scala 111:{38,38}]
  wire  _GEN_743 = 7'h60 == reqIndex ? way1Age_96 : _GEN_742; // @[ICache.scala 111:{38,38}]
  wire  _GEN_744 = 7'h61 == reqIndex ? way1Age_97 : _GEN_743; // @[ICache.scala 111:{38,38}]
  wire  _GEN_745 = 7'h62 == reqIndex ? way1Age_98 : _GEN_744; // @[ICache.scala 111:{38,38}]
  wire  _GEN_746 = 7'h63 == reqIndex ? way1Age_99 : _GEN_745; // @[ICache.scala 111:{38,38}]
  wire  _GEN_747 = 7'h64 == reqIndex ? way1Age_100 : _GEN_746; // @[ICache.scala 111:{38,38}]
  wire  _GEN_748 = 7'h65 == reqIndex ? way1Age_101 : _GEN_747; // @[ICache.scala 111:{38,38}]
  wire  _GEN_749 = 7'h66 == reqIndex ? way1Age_102 : _GEN_748; // @[ICache.scala 111:{38,38}]
  wire  _GEN_750 = 7'h67 == reqIndex ? way1Age_103 : _GEN_749; // @[ICache.scala 111:{38,38}]
  wire  _GEN_751 = 7'h68 == reqIndex ? way1Age_104 : _GEN_750; // @[ICache.scala 111:{38,38}]
  wire  _GEN_752 = 7'h69 == reqIndex ? way1Age_105 : _GEN_751; // @[ICache.scala 111:{38,38}]
  wire  _GEN_753 = 7'h6a == reqIndex ? way1Age_106 : _GEN_752; // @[ICache.scala 111:{38,38}]
  wire  _GEN_754 = 7'h6b == reqIndex ? way1Age_107 : _GEN_753; // @[ICache.scala 111:{38,38}]
  wire  _GEN_755 = 7'h6c == reqIndex ? way1Age_108 : _GEN_754; // @[ICache.scala 111:{38,38}]
  wire  _GEN_756 = 7'h6d == reqIndex ? way1Age_109 : _GEN_755; // @[ICache.scala 111:{38,38}]
  wire  _GEN_757 = 7'h6e == reqIndex ? way1Age_110 : _GEN_756; // @[ICache.scala 111:{38,38}]
  wire  _GEN_758 = 7'h6f == reqIndex ? way1Age_111 : _GEN_757; // @[ICache.scala 111:{38,38}]
  wire  _GEN_759 = 7'h70 == reqIndex ? way1Age_112 : _GEN_758; // @[ICache.scala 111:{38,38}]
  wire  _GEN_760 = 7'h71 == reqIndex ? way1Age_113 : _GEN_759; // @[ICache.scala 111:{38,38}]
  wire  _GEN_761 = 7'h72 == reqIndex ? way1Age_114 : _GEN_760; // @[ICache.scala 111:{38,38}]
  wire  _GEN_762 = 7'h73 == reqIndex ? way1Age_115 : _GEN_761; // @[ICache.scala 111:{38,38}]
  wire  _GEN_763 = 7'h74 == reqIndex ? way1Age_116 : _GEN_762; // @[ICache.scala 111:{38,38}]
  wire  _GEN_764 = 7'h75 == reqIndex ? way1Age_117 : _GEN_763; // @[ICache.scala 111:{38,38}]
  wire  _GEN_765 = 7'h76 == reqIndex ? way1Age_118 : _GEN_764; // @[ICache.scala 111:{38,38}]
  wire  _GEN_766 = 7'h77 == reqIndex ? way1Age_119 : _GEN_765; // @[ICache.scala 111:{38,38}]
  wire  _GEN_767 = 7'h78 == reqIndex ? way1Age_120 : _GEN_766; // @[ICache.scala 111:{38,38}]
  wire  _GEN_768 = 7'h79 == reqIndex ? way1Age_121 : _GEN_767; // @[ICache.scala 111:{38,38}]
  wire  _GEN_769 = 7'h7a == reqIndex ? way1Age_122 : _GEN_768; // @[ICache.scala 111:{38,38}]
  wire  _GEN_770 = 7'h7b == reqIndex ? way1Age_123 : _GEN_769; // @[ICache.scala 111:{38,38}]
  wire  _GEN_771 = 7'h7c == reqIndex ? way1Age_124 : _GEN_770; // @[ICache.scala 111:{38,38}]
  wire  _GEN_772 = 7'h7d == reqIndex ? way1Age_125 : _GEN_771; // @[ICache.scala 111:{38,38}]
  wire  _GEN_773 = 7'h7e == reqIndex ? way1Age_126 : _GEN_772; // @[ICache.scala 111:{38,38}]
  wire  _GEN_774 = 7'h7f == reqIndex ? way1Age_127 : _GEN_773; // @[ICache.scala 111:{38,38}]
  wire  ageWay1En = ~_GEN_774 & sFillEn; // @[ICache.scala 111:47]
  wire  _GEN_2311 = 7'h0 == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1159 = 7'h0 == reqIndex | way0V_0; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2312 = 7'h1 == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1160 = 7'h1 == reqIndex | way0V_1; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2313 = 7'h2 == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1161 = 7'h2 == reqIndex | way0V_2; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2314 = 7'h3 == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1162 = 7'h3 == reqIndex | way0V_3; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2315 = 7'h4 == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1163 = 7'h4 == reqIndex | way0V_4; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2316 = 7'h5 == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1164 = 7'h5 == reqIndex | way0V_5; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2317 = 7'h6 == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1165 = 7'h6 == reqIndex | way0V_6; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2318 = 7'h7 == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1166 = 7'h7 == reqIndex | way0V_7; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2319 = 7'h8 == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1167 = 7'h8 == reqIndex | way0V_8; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2320 = 7'h9 == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1168 = 7'h9 == reqIndex | way0V_9; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2321 = 7'ha == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1169 = 7'ha == reqIndex | way0V_10; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2322 = 7'hb == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1170 = 7'hb == reqIndex | way0V_11; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2323 = 7'hc == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1171 = 7'hc == reqIndex | way0V_12; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2324 = 7'hd == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1172 = 7'hd == reqIndex | way0V_13; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2325 = 7'he == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1173 = 7'he == reqIndex | way0V_14; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2326 = 7'hf == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1174 = 7'hf == reqIndex | way0V_15; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2327 = 7'h10 == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1175 = 7'h10 == reqIndex | way0V_16; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2328 = 7'h11 == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1176 = 7'h11 == reqIndex | way0V_17; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2329 = 7'h12 == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1177 = 7'h12 == reqIndex | way0V_18; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2330 = 7'h13 == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1178 = 7'h13 == reqIndex | way0V_19; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2331 = 7'h14 == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1179 = 7'h14 == reqIndex | way0V_20; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2332 = 7'h15 == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1180 = 7'h15 == reqIndex | way0V_21; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2333 = 7'h16 == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1181 = 7'h16 == reqIndex | way0V_22; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2334 = 7'h17 == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1182 = 7'h17 == reqIndex | way0V_23; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2335 = 7'h18 == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1183 = 7'h18 == reqIndex | way0V_24; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2336 = 7'h19 == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1184 = 7'h19 == reqIndex | way0V_25; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2337 = 7'h1a == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1185 = 7'h1a == reqIndex | way0V_26; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2338 = 7'h1b == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1186 = 7'h1b == reqIndex | way0V_27; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2339 = 7'h1c == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1187 = 7'h1c == reqIndex | way0V_28; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2340 = 7'h1d == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1188 = 7'h1d == reqIndex | way0V_29; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2341 = 7'h1e == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1189 = 7'h1e == reqIndex | way0V_30; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2342 = 7'h1f == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1190 = 7'h1f == reqIndex | way0V_31; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2343 = 7'h20 == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1191 = 7'h20 == reqIndex | way0V_32; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2344 = 7'h21 == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1192 = 7'h21 == reqIndex | way0V_33; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2345 = 7'h22 == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1193 = 7'h22 == reqIndex | way0V_34; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2346 = 7'h23 == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1194 = 7'h23 == reqIndex | way0V_35; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2347 = 7'h24 == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1195 = 7'h24 == reqIndex | way0V_36; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2348 = 7'h25 == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1196 = 7'h25 == reqIndex | way0V_37; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2349 = 7'h26 == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1197 = 7'h26 == reqIndex | way0V_38; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2350 = 7'h27 == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1198 = 7'h27 == reqIndex | way0V_39; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2351 = 7'h28 == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1199 = 7'h28 == reqIndex | way0V_40; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2352 = 7'h29 == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1200 = 7'h29 == reqIndex | way0V_41; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2353 = 7'h2a == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1201 = 7'h2a == reqIndex | way0V_42; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2354 = 7'h2b == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1202 = 7'h2b == reqIndex | way0V_43; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2355 = 7'h2c == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1203 = 7'h2c == reqIndex | way0V_44; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2356 = 7'h2d == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1204 = 7'h2d == reqIndex | way0V_45; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2357 = 7'h2e == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1205 = 7'h2e == reqIndex | way0V_46; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2358 = 7'h2f == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1206 = 7'h2f == reqIndex | way0V_47; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2359 = 7'h30 == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1207 = 7'h30 == reqIndex | way0V_48; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2360 = 7'h31 == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1208 = 7'h31 == reqIndex | way0V_49; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2361 = 7'h32 == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1209 = 7'h32 == reqIndex | way0V_50; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2362 = 7'h33 == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1210 = 7'h33 == reqIndex | way0V_51; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2363 = 7'h34 == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1211 = 7'h34 == reqIndex | way0V_52; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2364 = 7'h35 == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1212 = 7'h35 == reqIndex | way0V_53; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2365 = 7'h36 == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1213 = 7'h36 == reqIndex | way0V_54; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2366 = 7'h37 == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1214 = 7'h37 == reqIndex | way0V_55; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2367 = 7'h38 == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1215 = 7'h38 == reqIndex | way0V_56; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2368 = 7'h39 == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1216 = 7'h39 == reqIndex | way0V_57; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2369 = 7'h3a == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1217 = 7'h3a == reqIndex | way0V_58; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2370 = 7'h3b == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1218 = 7'h3b == reqIndex | way0V_59; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2371 = 7'h3c == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1219 = 7'h3c == reqIndex | way0V_60; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2372 = 7'h3d == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1220 = 7'h3d == reqIndex | way0V_61; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2373 = 7'h3e == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1221 = 7'h3e == reqIndex | way0V_62; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2374 = 7'h3f == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1222 = 7'h3f == reqIndex | way0V_63; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2375 = 7'h40 == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1223 = 7'h40 == reqIndex | way0V_64; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2376 = 7'h41 == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1224 = 7'h41 == reqIndex | way0V_65; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2377 = 7'h42 == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1225 = 7'h42 == reqIndex | way0V_66; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2378 = 7'h43 == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1226 = 7'h43 == reqIndex | way0V_67; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2379 = 7'h44 == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1227 = 7'h44 == reqIndex | way0V_68; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2380 = 7'h45 == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1228 = 7'h45 == reqIndex | way0V_69; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2381 = 7'h46 == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1229 = 7'h46 == reqIndex | way0V_70; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2382 = 7'h47 == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1230 = 7'h47 == reqIndex | way0V_71; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2383 = 7'h48 == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1231 = 7'h48 == reqIndex | way0V_72; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2384 = 7'h49 == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1232 = 7'h49 == reqIndex | way0V_73; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2385 = 7'h4a == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1233 = 7'h4a == reqIndex | way0V_74; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2386 = 7'h4b == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1234 = 7'h4b == reqIndex | way0V_75; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2387 = 7'h4c == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1235 = 7'h4c == reqIndex | way0V_76; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2388 = 7'h4d == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1236 = 7'h4d == reqIndex | way0V_77; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2389 = 7'h4e == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1237 = 7'h4e == reqIndex | way0V_78; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2390 = 7'h4f == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1238 = 7'h4f == reqIndex | way0V_79; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2391 = 7'h50 == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1239 = 7'h50 == reqIndex | way0V_80; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2392 = 7'h51 == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1240 = 7'h51 == reqIndex | way0V_81; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2393 = 7'h52 == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1241 = 7'h52 == reqIndex | way0V_82; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2394 = 7'h53 == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1242 = 7'h53 == reqIndex | way0V_83; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2395 = 7'h54 == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1243 = 7'h54 == reqIndex | way0V_84; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2396 = 7'h55 == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1244 = 7'h55 == reqIndex | way0V_85; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2397 = 7'h56 == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1245 = 7'h56 == reqIndex | way0V_86; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2398 = 7'h57 == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1246 = 7'h57 == reqIndex | way0V_87; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2399 = 7'h58 == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1247 = 7'h58 == reqIndex | way0V_88; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2400 = 7'h59 == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1248 = 7'h59 == reqIndex | way0V_89; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2401 = 7'h5a == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1249 = 7'h5a == reqIndex | way0V_90; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2402 = 7'h5b == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1250 = 7'h5b == reqIndex | way0V_91; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2403 = 7'h5c == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1251 = 7'h5c == reqIndex | way0V_92; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2404 = 7'h5d == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1252 = 7'h5d == reqIndex | way0V_93; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2405 = 7'h5e == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1253 = 7'h5e == reqIndex | way0V_94; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2406 = 7'h5f == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1254 = 7'h5f == reqIndex | way0V_95; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2407 = 7'h60 == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1255 = 7'h60 == reqIndex | way0V_96; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2408 = 7'h61 == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1256 = 7'h61 == reqIndex | way0V_97; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2409 = 7'h62 == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1257 = 7'h62 == reqIndex | way0V_98; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2410 = 7'h63 == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1258 = 7'h63 == reqIndex | way0V_99; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2411 = 7'h64 == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1259 = 7'h64 == reqIndex | way0V_100; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2412 = 7'h65 == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1260 = 7'h65 == reqIndex | way0V_101; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2413 = 7'h66 == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1261 = 7'h66 == reqIndex | way0V_102; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2414 = 7'h67 == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1262 = 7'h67 == reqIndex | way0V_103; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2415 = 7'h68 == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1263 = 7'h68 == reqIndex | way0V_104; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2416 = 7'h69 == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1264 = 7'h69 == reqIndex | way0V_105; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2417 = 7'h6a == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1265 = 7'h6a == reqIndex | way0V_106; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2418 = 7'h6b == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1266 = 7'h6b == reqIndex | way0V_107; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2419 = 7'h6c == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1267 = 7'h6c == reqIndex | way0V_108; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2420 = 7'h6d == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1268 = 7'h6d == reqIndex | way0V_109; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2421 = 7'h6e == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1269 = 7'h6e == reqIndex | way0V_110; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2422 = 7'h6f == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1270 = 7'h6f == reqIndex | way0V_111; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2423 = 7'h70 == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1271 = 7'h70 == reqIndex | way0V_112; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2424 = 7'h71 == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1272 = 7'h71 == reqIndex | way0V_113; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2425 = 7'h72 == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1273 = 7'h72 == reqIndex | way0V_114; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2426 = 7'h73 == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1274 = 7'h73 == reqIndex | way0V_115; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2427 = 7'h74 == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1275 = 7'h74 == reqIndex | way0V_116; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2428 = 7'h75 == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1276 = 7'h75 == reqIndex | way0V_117; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2429 = 7'h76 == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1277 = 7'h76 == reqIndex | way0V_118; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2430 = 7'h77 == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1278 = 7'h77 == reqIndex | way0V_119; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2431 = 7'h78 == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1279 = 7'h78 == reqIndex | way0V_120; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2432 = 7'h79 == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1280 = 7'h79 == reqIndex | way0V_121; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2433 = 7'h7a == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1281 = 7'h7a == reqIndex | way0V_122; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2434 = 7'h7b == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1282 = 7'h7b == reqIndex | way0V_123; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2435 = 7'h7c == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1283 = 7'h7c == reqIndex | way0V_124; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2436 = 7'h7d == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1284 = 7'h7d == reqIndex | way0V_125; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2437 = 7'h7e == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1285 = 7'h7e == reqIndex | way0V_126; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_2438 = 7'h7f == reqIndex; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1286 = 7'h7f == reqIndex | way0V_127; // @[ICache.scala 120:{21,21} 27:22]
  wire  _GEN_1415 = _GEN_2311 | way1V_0; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1416 = _GEN_2312 | way1V_1; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1417 = _GEN_2313 | way1V_2; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1418 = _GEN_2314 | way1V_3; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1419 = _GEN_2315 | way1V_4; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1420 = _GEN_2316 | way1V_5; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1421 = _GEN_2317 | way1V_6; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1422 = _GEN_2318 | way1V_7; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1423 = _GEN_2319 | way1V_8; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1424 = _GEN_2320 | way1V_9; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1425 = _GEN_2321 | way1V_10; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1426 = _GEN_2322 | way1V_11; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1427 = _GEN_2323 | way1V_12; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1428 = _GEN_2324 | way1V_13; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1429 = _GEN_2325 | way1V_14; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1430 = _GEN_2326 | way1V_15; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1431 = _GEN_2327 | way1V_16; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1432 = _GEN_2328 | way1V_17; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1433 = _GEN_2329 | way1V_18; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1434 = _GEN_2330 | way1V_19; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1435 = _GEN_2331 | way1V_20; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1436 = _GEN_2332 | way1V_21; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1437 = _GEN_2333 | way1V_22; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1438 = _GEN_2334 | way1V_23; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1439 = _GEN_2335 | way1V_24; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1440 = _GEN_2336 | way1V_25; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1441 = _GEN_2337 | way1V_26; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1442 = _GEN_2338 | way1V_27; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1443 = _GEN_2339 | way1V_28; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1444 = _GEN_2340 | way1V_29; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1445 = _GEN_2341 | way1V_30; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1446 = _GEN_2342 | way1V_31; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1447 = _GEN_2343 | way1V_32; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1448 = _GEN_2344 | way1V_33; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1449 = _GEN_2345 | way1V_34; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1450 = _GEN_2346 | way1V_35; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1451 = _GEN_2347 | way1V_36; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1452 = _GEN_2348 | way1V_37; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1453 = _GEN_2349 | way1V_38; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1454 = _GEN_2350 | way1V_39; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1455 = _GEN_2351 | way1V_40; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1456 = _GEN_2352 | way1V_41; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1457 = _GEN_2353 | way1V_42; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1458 = _GEN_2354 | way1V_43; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1459 = _GEN_2355 | way1V_44; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1460 = _GEN_2356 | way1V_45; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1461 = _GEN_2357 | way1V_46; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1462 = _GEN_2358 | way1V_47; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1463 = _GEN_2359 | way1V_48; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1464 = _GEN_2360 | way1V_49; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1465 = _GEN_2361 | way1V_50; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1466 = _GEN_2362 | way1V_51; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1467 = _GEN_2363 | way1V_52; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1468 = _GEN_2364 | way1V_53; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1469 = _GEN_2365 | way1V_54; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1470 = _GEN_2366 | way1V_55; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1471 = _GEN_2367 | way1V_56; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1472 = _GEN_2368 | way1V_57; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1473 = _GEN_2369 | way1V_58; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1474 = _GEN_2370 | way1V_59; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1475 = _GEN_2371 | way1V_60; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1476 = _GEN_2372 | way1V_61; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1477 = _GEN_2373 | way1V_62; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1478 = _GEN_2374 | way1V_63; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1479 = _GEN_2375 | way1V_64; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1480 = _GEN_2376 | way1V_65; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1481 = _GEN_2377 | way1V_66; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1482 = _GEN_2378 | way1V_67; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1483 = _GEN_2379 | way1V_68; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1484 = _GEN_2380 | way1V_69; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1485 = _GEN_2381 | way1V_70; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1486 = _GEN_2382 | way1V_71; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1487 = _GEN_2383 | way1V_72; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1488 = _GEN_2384 | way1V_73; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1489 = _GEN_2385 | way1V_74; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1490 = _GEN_2386 | way1V_75; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1491 = _GEN_2387 | way1V_76; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1492 = _GEN_2388 | way1V_77; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1493 = _GEN_2389 | way1V_78; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1494 = _GEN_2390 | way1V_79; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1495 = _GEN_2391 | way1V_80; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1496 = _GEN_2392 | way1V_81; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1497 = _GEN_2393 | way1V_82; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1498 = _GEN_2394 | way1V_83; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1499 = _GEN_2395 | way1V_84; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1500 = _GEN_2396 | way1V_85; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1501 = _GEN_2397 | way1V_86; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1502 = _GEN_2398 | way1V_87; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1503 = _GEN_2399 | way1V_88; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1504 = _GEN_2400 | way1V_89; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1505 = _GEN_2401 | way1V_90; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1506 = _GEN_2402 | way1V_91; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1507 = _GEN_2403 | way1V_92; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1508 = _GEN_2404 | way1V_93; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1509 = _GEN_2405 | way1V_94; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1510 = _GEN_2406 | way1V_95; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1511 = _GEN_2407 | way1V_96; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1512 = _GEN_2408 | way1V_97; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1513 = _GEN_2409 | way1V_98; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1514 = _GEN_2410 | way1V_99; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1515 = _GEN_2411 | way1V_100; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1516 = _GEN_2412 | way1V_101; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1517 = _GEN_2413 | way1V_102; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1518 = _GEN_2414 | way1V_103; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1519 = _GEN_2415 | way1V_104; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1520 = _GEN_2416 | way1V_105; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1521 = _GEN_2417 | way1V_106; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1522 = _GEN_2418 | way1V_107; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1523 = _GEN_2419 | way1V_108; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1524 = _GEN_2420 | way1V_109; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1525 = _GEN_2421 | way1V_110; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1526 = _GEN_2422 | way1V_111; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1527 = _GEN_2423 | way1V_112; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1528 = _GEN_2424 | way1V_113; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1529 = _GEN_2425 | way1V_114; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1530 = _GEN_2426 | way1V_115; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1531 = _GEN_2427 | way1V_116; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1532 = _GEN_2428 | way1V_117; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1533 = _GEN_2429 | way1V_118; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1534 = _GEN_2430 | way1V_119; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1535 = _GEN_2431 | way1V_120; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1536 = _GEN_2432 | way1V_121; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1537 = _GEN_2433 | way1V_122; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1538 = _GEN_2434 | way1V_123; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1539 = _GEN_2435 | way1V_124; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1540 = _GEN_2436 | way1V_125; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1541 = _GEN_2437 | way1V_126; // @[ICache.scala 123:{21,21} 32:22]
  wire  _GEN_1542 = _GEN_2438 | way1V_127; // @[ICache.scala 123:{21,21} 32:22]
  S011HD1P_X32Y2D128 req ( // @[ICache.scala 54:19]
    .Q(req_Q),
    .CLK(req_CLK),
    .CEN(req_CEN),
    .WEN(req_WEN),
    .A(req_A),
    .D(req_D)
  );
  assign io_imem_inst_ready = sReadEn & cacheHitEn; // @[ICache.scala 92:28]
  assign io_imem_inst_read = 2'h3 == reqOff[3:2] ? rData[127:96] : _io_imem_inst_read_T_8; // @[Mux.scala 81:58]
  assign io_out_inst_valid = state == 2'h2; // @[ICache.scala 100:22]
  assign io_out_inst_addr = sAxiEn ? io_imem_inst_addr : 32'h0; // @[ICache.scala 103:23]
  assign req_CLK = clock; // @[ICache.scala 55:14]
  assign req_CEN = 1'h1; // @[ICache.scala 56:14]
  assign req_WEN = state == 2'h3; // @[ICache.scala 108:23]
  assign req_A = ~sFillEn ? cacheRIndex : cacheWIndex; // @[ICache.scala 58:20]
  assign req_D = cacheWData; // @[ICache.scala 59:14]
  always @(posedge clock) begin
    if (reset) begin // @[ICache.scala 22:27]
      cacheWData <= 128'h0; // @[ICache.scala 22:27]
    end else if (sAxiEn & io_out_inst_ready) begin // @[ICache.scala 105:20]
      cacheWData <= io_out_inst_read;
    end else begin
      cacheWData <= 128'h0;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_0 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_0 <= _GEN_1159;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_1 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_1 <= _GEN_1160;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_2 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_2 <= _GEN_1161;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_3 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_3 <= _GEN_1162;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_4 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_4 <= _GEN_1163;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_5 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_5 <= _GEN_1164;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_6 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_6 <= _GEN_1165;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_7 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_7 <= _GEN_1166;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_8 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_8 <= _GEN_1167;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_9 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_9 <= _GEN_1168;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_10 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_10 <= _GEN_1169;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_11 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_11 <= _GEN_1170;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_12 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_12 <= _GEN_1171;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_13 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_13 <= _GEN_1172;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_14 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_14 <= _GEN_1173;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_15 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_15 <= _GEN_1174;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_16 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_16 <= _GEN_1175;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_17 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_17 <= _GEN_1176;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_18 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_18 <= _GEN_1177;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_19 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_19 <= _GEN_1178;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_20 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_20 <= _GEN_1179;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_21 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_21 <= _GEN_1180;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_22 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_22 <= _GEN_1181;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_23 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_23 <= _GEN_1182;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_24 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_24 <= _GEN_1183;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_25 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_25 <= _GEN_1184;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_26 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_26 <= _GEN_1185;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_27 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_27 <= _GEN_1186;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_28 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_28 <= _GEN_1187;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_29 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_29 <= _GEN_1188;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_30 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_30 <= _GEN_1189;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_31 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_31 <= _GEN_1190;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_32 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_32 <= _GEN_1191;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_33 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_33 <= _GEN_1192;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_34 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_34 <= _GEN_1193;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_35 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_35 <= _GEN_1194;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_36 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_36 <= _GEN_1195;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_37 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_37 <= _GEN_1196;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_38 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_38 <= _GEN_1197;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_39 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_39 <= _GEN_1198;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_40 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_40 <= _GEN_1199;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_41 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_41 <= _GEN_1200;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_42 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_42 <= _GEN_1201;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_43 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_43 <= _GEN_1202;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_44 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_44 <= _GEN_1203;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_45 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_45 <= _GEN_1204;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_46 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_46 <= _GEN_1205;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_47 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_47 <= _GEN_1206;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_48 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_48 <= _GEN_1207;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_49 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_49 <= _GEN_1208;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_50 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_50 <= _GEN_1209;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_51 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_51 <= _GEN_1210;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_52 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_52 <= _GEN_1211;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_53 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_53 <= _GEN_1212;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_54 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_54 <= _GEN_1213;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_55 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_55 <= _GEN_1214;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_56 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_56 <= _GEN_1215;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_57 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_57 <= _GEN_1216;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_58 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_58 <= _GEN_1217;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_59 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_59 <= _GEN_1218;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_60 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_60 <= _GEN_1219;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_61 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_61 <= _GEN_1220;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_62 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_62 <= _GEN_1221;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_63 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_63 <= _GEN_1222;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_64 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_64 <= _GEN_1223;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_65 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_65 <= _GEN_1224;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_66 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_66 <= _GEN_1225;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_67 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_67 <= _GEN_1226;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_68 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_68 <= _GEN_1227;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_69 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_69 <= _GEN_1228;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_70 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_70 <= _GEN_1229;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_71 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_71 <= _GEN_1230;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_72 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_72 <= _GEN_1231;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_73 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_73 <= _GEN_1232;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_74 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_74 <= _GEN_1233;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_75 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_75 <= _GEN_1234;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_76 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_76 <= _GEN_1235;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_77 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_77 <= _GEN_1236;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_78 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_78 <= _GEN_1237;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_79 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_79 <= _GEN_1238;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_80 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_80 <= _GEN_1239;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_81 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_81 <= _GEN_1240;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_82 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_82 <= _GEN_1241;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_83 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_83 <= _GEN_1242;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_84 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_84 <= _GEN_1243;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_85 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_85 <= _GEN_1244;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_86 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_86 <= _GEN_1245;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_87 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_87 <= _GEN_1246;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_88 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_88 <= _GEN_1247;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_89 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_89 <= _GEN_1248;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_90 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_90 <= _GEN_1249;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_91 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_91 <= _GEN_1250;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_92 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_92 <= _GEN_1251;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_93 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_93 <= _GEN_1252;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_94 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_94 <= _GEN_1253;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_95 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_95 <= _GEN_1254;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_96 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_96 <= _GEN_1255;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_97 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_97 <= _GEN_1256;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_98 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_98 <= _GEN_1257;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_99 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_99 <= _GEN_1258;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_100 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_100 <= _GEN_1259;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_101 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_101 <= _GEN_1260;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_102 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_102 <= _GEN_1261;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_103 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_103 <= _GEN_1262;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_104 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_104 <= _GEN_1263;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_105 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_105 <= _GEN_1264;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_106 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_106 <= _GEN_1265;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_107 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_107 <= _GEN_1266;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_108 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_108 <= _GEN_1267;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_109 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_109 <= _GEN_1268;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_110 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_110 <= _GEN_1269;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_111 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_111 <= _GEN_1270;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_112 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_112 <= _GEN_1271;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_113 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_113 <= _GEN_1272;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_114 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_114 <= _GEN_1273;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_115 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_115 <= _GEN_1274;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_116 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_116 <= _GEN_1275;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_117 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_117 <= _GEN_1276;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_118 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_118 <= _GEN_1277;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_119 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_119 <= _GEN_1278;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_120 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_120 <= _GEN_1279;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_121 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_121 <= _GEN_1280;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_122 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_122 <= _GEN_1281;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_123 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_123 <= _GEN_1282;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_124 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_124 <= _GEN_1283;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_125 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_125 <= _GEN_1284;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_126 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_126 <= _GEN_1285;
    end
    if (reset) begin // @[ICache.scala 27:22]
      way0V_127 <= 1'h0; // @[ICache.scala 27:22]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      way0V_127 <= _GEN_1286;
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_0 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h0 == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_0 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_1 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h1 == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_1 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_2 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h2 == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_2 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_3 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h3 == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_3 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_4 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h4 == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_4 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_5 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h5 == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_5 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_6 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h6 == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_6 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_7 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h7 == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_7 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_8 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h8 == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_8 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_9 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h9 == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_9 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_10 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'ha == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_10 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_11 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'hb == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_11 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_12 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'hc == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_12 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_13 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'hd == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_13 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_14 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'he == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_14 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_15 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'hf == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_15 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_16 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h10 == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_16 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_17 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h11 == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_17 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_18 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h12 == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_18 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_19 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h13 == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_19 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_20 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h14 == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_20 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_21 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h15 == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_21 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_22 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h16 == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_22 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_23 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h17 == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_23 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_24 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h18 == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_24 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_25 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h19 == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_25 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_26 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h1a == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_26 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_27 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h1b == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_27 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_28 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h1c == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_28 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_29 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h1d == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_29 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_30 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h1e == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_30 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_31 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h1f == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_31 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_32 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h20 == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_32 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_33 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h21 == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_33 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_34 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h22 == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_34 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_35 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h23 == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_35 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_36 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h24 == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_36 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_37 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h25 == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_37 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_38 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h26 == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_38 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_39 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h27 == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_39 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_40 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h28 == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_40 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_41 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h29 == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_41 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_42 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h2a == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_42 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_43 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h2b == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_43 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_44 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h2c == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_44 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_45 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h2d == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_45 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_46 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h2e == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_46 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_47 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h2f == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_47 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_48 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h30 == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_48 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_49 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h31 == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_49 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_50 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h32 == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_50 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_51 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h33 == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_51 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_52 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h34 == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_52 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_53 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h35 == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_53 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_54 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h36 == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_54 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_55 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h37 == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_55 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_56 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h38 == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_56 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_57 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h39 == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_57 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_58 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h3a == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_58 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_59 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h3b == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_59 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_60 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h3c == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_60 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_61 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h3d == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_61 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_62 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h3e == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_62 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_63 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h3f == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_63 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_64 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h40 == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_64 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_65 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h41 == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_65 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_66 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h42 == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_66 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_67 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h43 == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_67 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_68 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h44 == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_68 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_69 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h45 == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_69 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_70 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h46 == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_70 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_71 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h47 == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_71 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_72 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h48 == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_72 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_73 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h49 == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_73 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_74 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h4a == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_74 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_75 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h4b == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_75 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_76 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h4c == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_76 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_77 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h4d == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_77 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_78 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h4e == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_78 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_79 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h4f == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_79 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_80 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h50 == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_80 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_81 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h51 == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_81 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_82 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h52 == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_82 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_83 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h53 == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_83 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_84 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h54 == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_84 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_85 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h55 == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_85 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_86 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h56 == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_86 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_87 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h57 == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_87 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_88 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h58 == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_88 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_89 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h59 == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_89 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_90 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h5a == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_90 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_91 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h5b == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_91 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_92 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h5c == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_92 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_93 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h5d == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_93 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_94 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h5e == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_94 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_95 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h5f == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_95 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_96 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h60 == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_96 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_97 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h61 == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_97 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_98 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h62 == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_98 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_99 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h63 == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_99 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_100 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h64 == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_100 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_101 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h65 == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_101 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_102 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h66 == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_102 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_103 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h67 == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_103 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_104 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h68 == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_104 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_105 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h69 == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_105 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_106 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h6a == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_106 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_107 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h6b == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_107 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_108 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h6c == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_108 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_109 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h6d == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_109 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_110 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h6e == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_110 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_111 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h6f == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_111 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_112 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h70 == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_112 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_113 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h71 == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_113 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_114 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h72 == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_114 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_115 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h73 == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_115 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_116 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h74 == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_116 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_117 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h75 == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_117 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_118 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h76 == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_118 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_119 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h77 == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_119 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_120 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h78 == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_120 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_121 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h79 == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_121 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_122 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h7a == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_122 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_123 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h7b == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_123 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_124 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h7c == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_124 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_125 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h7d == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_125 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_126 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h7e == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_126 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 28:24]
      way0Tag_127 <= 21'h0; // @[ICache.scala 28:24]
    end else if (ageWay0En) begin // @[ICache.scala 118:19]
      if (7'h7f == reqIndex) begin // @[ICache.scala 119:23]
        way0Tag_127 <= reqTag; // @[ICache.scala 119:23]
      end
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_0 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h0 == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_0 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_1 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h1 == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_1 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_2 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h2 == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_2 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_3 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h3 == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_3 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_4 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h4 == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_4 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_5 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h5 == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_5 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_6 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h6 == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_6 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_7 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h7 == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_7 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_8 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h8 == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_8 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_9 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h9 == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_9 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_10 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'ha == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_10 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_11 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'hb == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_11 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_12 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'hc == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_12 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_13 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'hd == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_13 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_14 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'he == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_14 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_15 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'hf == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_15 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_16 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h10 == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_16 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_17 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h11 == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_17 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_18 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h12 == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_18 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_19 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h13 == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_19 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_20 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h14 == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_20 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_21 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h15 == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_21 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_22 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h16 == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_22 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_23 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h17 == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_23 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_24 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h18 == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_24 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_25 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h19 == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_25 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_26 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h1a == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_26 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_27 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h1b == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_27 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_28 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h1c == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_28 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_29 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h1d == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_29 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_30 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h1e == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_30 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_31 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h1f == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_31 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_32 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h20 == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_32 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_33 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h21 == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_33 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_34 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h22 == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_34 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_35 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h23 == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_35 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_36 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h24 == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_36 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_37 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h25 == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_37 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_38 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h26 == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_38 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_39 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h27 == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_39 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_40 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h28 == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_40 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_41 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h29 == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_41 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_42 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h2a == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_42 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_43 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h2b == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_43 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_44 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h2c == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_44 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_45 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h2d == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_45 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_46 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h2e == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_46 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_47 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h2f == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_47 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_48 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h30 == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_48 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_49 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h31 == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_49 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_50 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h32 == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_50 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_51 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h33 == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_51 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_52 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h34 == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_52 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_53 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h35 == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_53 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_54 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h36 == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_54 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_55 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h37 == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_55 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_56 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h38 == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_56 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_57 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h39 == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_57 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_58 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h3a == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_58 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_59 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h3b == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_59 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_60 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h3c == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_60 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_61 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h3d == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_61 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_62 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h3e == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_62 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_63 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h3f == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_63 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_64 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h40 == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_64 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_65 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h41 == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_65 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_66 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h42 == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_66 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_67 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h43 == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_67 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_68 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h44 == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_68 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_69 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h45 == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_69 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_70 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h46 == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_70 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_71 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h47 == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_71 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_72 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h48 == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_72 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_73 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h49 == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_73 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_74 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h4a == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_74 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_75 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h4b == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_75 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_76 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h4c == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_76 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_77 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h4d == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_77 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_78 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h4e == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_78 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_79 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h4f == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_79 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_80 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h50 == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_80 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_81 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h51 == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_81 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_82 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h52 == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_82 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_83 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h53 == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_83 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_84 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h54 == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_84 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_85 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h55 == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_85 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_86 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h56 == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_86 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_87 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h57 == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_87 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_88 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h58 == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_88 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_89 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h59 == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_89 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_90 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h5a == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_90 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_91 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h5b == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_91 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_92 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h5c == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_92 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_93 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h5d == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_93 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_94 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h5e == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_94 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_95 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h5f == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_95 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_96 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h60 == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_96 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_97 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h61 == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_97 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_98 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h62 == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_98 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_99 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h63 == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_99 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_100 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h64 == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_100 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_101 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h65 == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_101 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_102 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h66 == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_102 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_103 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h67 == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_103 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_104 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h68 == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_104 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_105 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h69 == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_105 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_106 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h6a == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_106 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_107 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h6b == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_107 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_108 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h6c == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_108 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_109 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h6d == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_109 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_110 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h6e == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_110 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_111 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h6f == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_111 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_112 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h70 == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_112 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_113 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h71 == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_113 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_114 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h72 == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_114 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_115 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h73 == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_115 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_116 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h74 == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_116 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_117 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h75 == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_117 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_118 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h76 == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_118 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_119 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h77 == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_119 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_120 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h78 == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_120 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_121 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h79 == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_121 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_122 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h7a == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_122 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_123 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h7b == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_123 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_124 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h7c == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_124 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_125 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h7d == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_125 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_126 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h7e == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_126 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 30:24]
      way0Age_127 <= 1'h0; // @[ICache.scala 30:24]
    end else if (7'h7f == reqIndex) begin // @[ICache.scala 113:21]
      way0Age_127 <= ageWay0En; // @[ICache.scala 113:21]
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_0 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_0 <= _GEN_1415;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_1 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_1 <= _GEN_1416;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_2 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_2 <= _GEN_1417;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_3 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_3 <= _GEN_1418;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_4 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_4 <= _GEN_1419;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_5 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_5 <= _GEN_1420;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_6 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_6 <= _GEN_1421;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_7 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_7 <= _GEN_1422;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_8 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_8 <= _GEN_1423;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_9 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_9 <= _GEN_1424;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_10 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_10 <= _GEN_1425;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_11 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_11 <= _GEN_1426;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_12 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_12 <= _GEN_1427;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_13 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_13 <= _GEN_1428;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_14 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_14 <= _GEN_1429;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_15 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_15 <= _GEN_1430;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_16 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_16 <= _GEN_1431;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_17 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_17 <= _GEN_1432;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_18 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_18 <= _GEN_1433;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_19 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_19 <= _GEN_1434;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_20 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_20 <= _GEN_1435;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_21 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_21 <= _GEN_1436;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_22 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_22 <= _GEN_1437;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_23 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_23 <= _GEN_1438;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_24 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_24 <= _GEN_1439;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_25 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_25 <= _GEN_1440;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_26 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_26 <= _GEN_1441;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_27 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_27 <= _GEN_1442;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_28 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_28 <= _GEN_1443;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_29 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_29 <= _GEN_1444;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_30 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_30 <= _GEN_1445;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_31 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_31 <= _GEN_1446;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_32 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_32 <= _GEN_1447;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_33 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_33 <= _GEN_1448;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_34 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_34 <= _GEN_1449;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_35 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_35 <= _GEN_1450;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_36 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_36 <= _GEN_1451;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_37 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_37 <= _GEN_1452;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_38 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_38 <= _GEN_1453;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_39 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_39 <= _GEN_1454;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_40 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_40 <= _GEN_1455;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_41 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_41 <= _GEN_1456;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_42 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_42 <= _GEN_1457;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_43 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_43 <= _GEN_1458;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_44 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_44 <= _GEN_1459;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_45 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_45 <= _GEN_1460;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_46 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_46 <= _GEN_1461;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_47 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_47 <= _GEN_1462;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_48 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_48 <= _GEN_1463;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_49 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_49 <= _GEN_1464;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_50 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_50 <= _GEN_1465;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_51 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_51 <= _GEN_1466;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_52 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_52 <= _GEN_1467;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_53 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_53 <= _GEN_1468;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_54 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_54 <= _GEN_1469;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_55 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_55 <= _GEN_1470;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_56 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_56 <= _GEN_1471;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_57 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_57 <= _GEN_1472;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_58 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_58 <= _GEN_1473;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_59 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_59 <= _GEN_1474;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_60 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_60 <= _GEN_1475;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_61 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_61 <= _GEN_1476;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_62 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_62 <= _GEN_1477;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_63 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_63 <= _GEN_1478;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_64 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_64 <= _GEN_1479;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_65 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_65 <= _GEN_1480;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_66 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_66 <= _GEN_1481;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_67 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_67 <= _GEN_1482;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_68 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_68 <= _GEN_1483;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_69 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_69 <= _GEN_1484;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_70 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_70 <= _GEN_1485;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_71 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_71 <= _GEN_1486;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_72 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_72 <= _GEN_1487;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_73 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_73 <= _GEN_1488;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_74 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_74 <= _GEN_1489;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_75 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_75 <= _GEN_1490;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_76 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_76 <= _GEN_1491;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_77 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_77 <= _GEN_1492;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_78 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_78 <= _GEN_1493;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_79 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_79 <= _GEN_1494;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_80 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_80 <= _GEN_1495;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_81 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_81 <= _GEN_1496;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_82 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_82 <= _GEN_1497;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_83 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_83 <= _GEN_1498;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_84 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_84 <= _GEN_1499;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_85 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_85 <= _GEN_1500;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_86 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_86 <= _GEN_1501;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_87 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_87 <= _GEN_1502;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_88 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_88 <= _GEN_1503;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_89 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_89 <= _GEN_1504;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_90 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_90 <= _GEN_1505;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_91 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_91 <= _GEN_1506;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_92 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_92 <= _GEN_1507;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_93 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_93 <= _GEN_1508;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_94 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_94 <= _GEN_1509;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_95 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_95 <= _GEN_1510;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_96 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_96 <= _GEN_1511;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_97 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_97 <= _GEN_1512;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_98 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_98 <= _GEN_1513;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_99 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_99 <= _GEN_1514;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_100 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_100 <= _GEN_1515;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_101 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_101 <= _GEN_1516;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_102 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_102 <= _GEN_1517;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_103 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_103 <= _GEN_1518;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_104 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_104 <= _GEN_1519;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_105 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_105 <= _GEN_1520;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_106 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_106 <= _GEN_1521;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_107 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_107 <= _GEN_1522;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_108 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_108 <= _GEN_1523;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_109 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_109 <= _GEN_1524;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_110 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_110 <= _GEN_1525;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_111 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_111 <= _GEN_1526;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_112 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_112 <= _GEN_1527;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_113 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_113 <= _GEN_1528;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_114 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_114 <= _GEN_1529;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_115 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_115 <= _GEN_1530;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_116 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_116 <= _GEN_1531;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_117 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_117 <= _GEN_1532;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_118 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_118 <= _GEN_1533;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_119 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_119 <= _GEN_1534;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_120 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_120 <= _GEN_1535;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_121 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_121 <= _GEN_1536;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_122 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_122 <= _GEN_1537;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_123 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_123 <= _GEN_1538;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_124 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_124 <= _GEN_1539;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_125 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_125 <= _GEN_1540;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_126 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_126 <= _GEN_1541;
      end
    end
    if (reset) begin // @[ICache.scala 32:22]
      way1V_127 <= 1'h0; // @[ICache.scala 32:22]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        way1V_127 <= _GEN_1542;
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_0 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h0 == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_0 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_1 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h1 == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_1 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_2 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h2 == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_2 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_3 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h3 == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_3 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_4 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h4 == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_4 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_5 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h5 == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_5 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_6 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h6 == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_6 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_7 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h7 == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_7 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_8 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h8 == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_8 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_9 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h9 == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_9 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_10 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'ha == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_10 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_11 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'hb == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_11 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_12 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'hc == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_12 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_13 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'hd == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_13 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_14 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'he == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_14 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_15 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'hf == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_15 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_16 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h10 == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_16 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_17 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h11 == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_17 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_18 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h12 == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_18 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_19 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h13 == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_19 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_20 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h14 == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_20 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_21 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h15 == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_21 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_22 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h16 == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_22 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_23 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h17 == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_23 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_24 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h18 == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_24 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_25 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h19 == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_25 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_26 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h1a == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_26 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_27 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h1b == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_27 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_28 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h1c == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_28 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_29 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h1d == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_29 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_30 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h1e == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_30 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_31 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h1f == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_31 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_32 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h20 == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_32 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_33 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h21 == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_33 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_34 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h22 == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_34 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_35 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h23 == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_35 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_36 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h24 == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_36 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_37 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h25 == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_37 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_38 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h26 == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_38 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_39 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h27 == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_39 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_40 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h28 == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_40 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_41 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h29 == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_41 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_42 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h2a == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_42 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_43 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h2b == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_43 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_44 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h2c == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_44 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_45 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h2d == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_45 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_46 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h2e == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_46 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_47 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h2f == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_47 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_48 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h30 == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_48 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_49 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h31 == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_49 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_50 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h32 == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_50 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_51 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h33 == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_51 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_52 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h34 == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_52 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_53 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h35 == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_53 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_54 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h36 == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_54 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_55 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h37 == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_55 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_56 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h38 == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_56 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_57 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h39 == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_57 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_58 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h3a == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_58 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_59 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h3b == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_59 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_60 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h3c == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_60 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_61 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h3d == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_61 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_62 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h3e == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_62 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_63 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h3f == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_63 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_64 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h40 == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_64 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_65 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h41 == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_65 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_66 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h42 == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_66 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_67 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h43 == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_67 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_68 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h44 == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_68 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_69 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h45 == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_69 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_70 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h46 == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_70 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_71 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h47 == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_71 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_72 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h48 == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_72 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_73 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h49 == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_73 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_74 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h4a == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_74 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_75 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h4b == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_75 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_76 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h4c == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_76 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_77 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h4d == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_77 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_78 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h4e == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_78 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_79 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h4f == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_79 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_80 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h50 == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_80 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_81 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h51 == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_81 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_82 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h52 == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_82 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_83 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h53 == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_83 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_84 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h54 == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_84 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_85 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h55 == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_85 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_86 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h56 == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_86 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_87 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h57 == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_87 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_88 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h58 == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_88 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_89 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h59 == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_89 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_90 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h5a == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_90 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_91 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h5b == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_91 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_92 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h5c == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_92 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_93 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h5d == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_93 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_94 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h5e == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_94 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_95 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h5f == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_95 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_96 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h60 == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_96 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_97 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h61 == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_97 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_98 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h62 == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_98 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_99 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h63 == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_99 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_100 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h64 == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_100 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_101 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h65 == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_101 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_102 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h66 == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_102 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_103 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h67 == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_103 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_104 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h68 == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_104 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_105 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h69 == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_105 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_106 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h6a == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_106 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_107 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h6b == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_107 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_108 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h6c == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_108 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_109 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h6d == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_109 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_110 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h6e == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_110 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_111 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h6f == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_111 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_112 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h70 == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_112 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_113 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h71 == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_113 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_114 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h72 == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_114 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_115 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h73 == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_115 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_116 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h74 == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_116 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_117 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h75 == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_117 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_118 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h76 == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_118 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_119 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h77 == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_119 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_120 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h78 == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_120 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_121 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h79 == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_121 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_122 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h7a == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_122 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_123 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h7b == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_123 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_124 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h7c == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_124 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_125 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h7d == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_125 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_126 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h7e == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_126 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 33:24]
      way1Tag_127 <= 21'h0; // @[ICache.scala 33:24]
    end else if (!(ageWay0En)) begin // @[ICache.scala 118:19]
      if (ageWay1En) begin // @[ICache.scala 121:26]
        if (7'h7f == reqIndex) begin // @[ICache.scala 122:23]
          way1Tag_127 <= reqTag; // @[ICache.scala 122:23]
        end
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_0 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h0 == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_0 <= 1'h0;
      end else begin
        way1Age_0 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_1 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h1 == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_1 <= 1'h0;
      end else begin
        way1Age_1 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_2 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h2 == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_2 <= 1'h0;
      end else begin
        way1Age_2 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_3 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h3 == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_3 <= 1'h0;
      end else begin
        way1Age_3 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_4 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h4 == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_4 <= 1'h0;
      end else begin
        way1Age_4 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_5 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h5 == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_5 <= 1'h0;
      end else begin
        way1Age_5 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_6 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h6 == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_6 <= 1'h0;
      end else begin
        way1Age_6 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_7 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h7 == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_7 <= 1'h0;
      end else begin
        way1Age_7 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_8 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h8 == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_8 <= 1'h0;
      end else begin
        way1Age_8 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_9 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h9 == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_9 <= 1'h0;
      end else begin
        way1Age_9 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_10 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'ha == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_10 <= 1'h0;
      end else begin
        way1Age_10 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_11 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'hb == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_11 <= 1'h0;
      end else begin
        way1Age_11 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_12 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'hc == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_12 <= 1'h0;
      end else begin
        way1Age_12 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_13 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'hd == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_13 <= 1'h0;
      end else begin
        way1Age_13 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_14 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'he == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_14 <= 1'h0;
      end else begin
        way1Age_14 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_15 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'hf == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_15 <= 1'h0;
      end else begin
        way1Age_15 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_16 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h10 == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_16 <= 1'h0;
      end else begin
        way1Age_16 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_17 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h11 == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_17 <= 1'h0;
      end else begin
        way1Age_17 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_18 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h12 == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_18 <= 1'h0;
      end else begin
        way1Age_18 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_19 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h13 == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_19 <= 1'h0;
      end else begin
        way1Age_19 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_20 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h14 == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_20 <= 1'h0;
      end else begin
        way1Age_20 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_21 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h15 == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_21 <= 1'h0;
      end else begin
        way1Age_21 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_22 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h16 == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_22 <= 1'h0;
      end else begin
        way1Age_22 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_23 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h17 == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_23 <= 1'h0;
      end else begin
        way1Age_23 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_24 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h18 == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_24 <= 1'h0;
      end else begin
        way1Age_24 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_25 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h19 == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_25 <= 1'h0;
      end else begin
        way1Age_25 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_26 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h1a == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_26 <= 1'h0;
      end else begin
        way1Age_26 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_27 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h1b == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_27 <= 1'h0;
      end else begin
        way1Age_27 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_28 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h1c == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_28 <= 1'h0;
      end else begin
        way1Age_28 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_29 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h1d == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_29 <= 1'h0;
      end else begin
        way1Age_29 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_30 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h1e == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_30 <= 1'h0;
      end else begin
        way1Age_30 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_31 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h1f == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_31 <= 1'h0;
      end else begin
        way1Age_31 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_32 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h20 == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_32 <= 1'h0;
      end else begin
        way1Age_32 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_33 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h21 == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_33 <= 1'h0;
      end else begin
        way1Age_33 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_34 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h22 == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_34 <= 1'h0;
      end else begin
        way1Age_34 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_35 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h23 == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_35 <= 1'h0;
      end else begin
        way1Age_35 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_36 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h24 == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_36 <= 1'h0;
      end else begin
        way1Age_36 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_37 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h25 == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_37 <= 1'h0;
      end else begin
        way1Age_37 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_38 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h26 == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_38 <= 1'h0;
      end else begin
        way1Age_38 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_39 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h27 == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_39 <= 1'h0;
      end else begin
        way1Age_39 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_40 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h28 == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_40 <= 1'h0;
      end else begin
        way1Age_40 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_41 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h29 == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_41 <= 1'h0;
      end else begin
        way1Age_41 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_42 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h2a == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_42 <= 1'h0;
      end else begin
        way1Age_42 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_43 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h2b == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_43 <= 1'h0;
      end else begin
        way1Age_43 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_44 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h2c == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_44 <= 1'h0;
      end else begin
        way1Age_44 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_45 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h2d == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_45 <= 1'h0;
      end else begin
        way1Age_45 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_46 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h2e == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_46 <= 1'h0;
      end else begin
        way1Age_46 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_47 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h2f == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_47 <= 1'h0;
      end else begin
        way1Age_47 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_48 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h30 == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_48 <= 1'h0;
      end else begin
        way1Age_48 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_49 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h31 == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_49 <= 1'h0;
      end else begin
        way1Age_49 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_50 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h32 == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_50 <= 1'h0;
      end else begin
        way1Age_50 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_51 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h33 == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_51 <= 1'h0;
      end else begin
        way1Age_51 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_52 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h34 == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_52 <= 1'h0;
      end else begin
        way1Age_52 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_53 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h35 == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_53 <= 1'h0;
      end else begin
        way1Age_53 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_54 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h36 == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_54 <= 1'h0;
      end else begin
        way1Age_54 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_55 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h37 == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_55 <= 1'h0;
      end else begin
        way1Age_55 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_56 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h38 == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_56 <= 1'h0;
      end else begin
        way1Age_56 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_57 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h39 == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_57 <= 1'h0;
      end else begin
        way1Age_57 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_58 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h3a == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_58 <= 1'h0;
      end else begin
        way1Age_58 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_59 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h3b == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_59 <= 1'h0;
      end else begin
        way1Age_59 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_60 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h3c == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_60 <= 1'h0;
      end else begin
        way1Age_60 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_61 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h3d == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_61 <= 1'h0;
      end else begin
        way1Age_61 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_62 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h3e == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_62 <= 1'h0;
      end else begin
        way1Age_62 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_63 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h3f == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_63 <= 1'h0;
      end else begin
        way1Age_63 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_64 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h40 == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_64 <= 1'h0;
      end else begin
        way1Age_64 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_65 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h41 == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_65 <= 1'h0;
      end else begin
        way1Age_65 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_66 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h42 == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_66 <= 1'h0;
      end else begin
        way1Age_66 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_67 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h43 == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_67 <= 1'h0;
      end else begin
        way1Age_67 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_68 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h44 == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_68 <= 1'h0;
      end else begin
        way1Age_68 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_69 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h45 == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_69 <= 1'h0;
      end else begin
        way1Age_69 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_70 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h46 == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_70 <= 1'h0;
      end else begin
        way1Age_70 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_71 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h47 == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_71 <= 1'h0;
      end else begin
        way1Age_71 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_72 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h48 == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_72 <= 1'h0;
      end else begin
        way1Age_72 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_73 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h49 == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_73 <= 1'h0;
      end else begin
        way1Age_73 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_74 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h4a == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_74 <= 1'h0;
      end else begin
        way1Age_74 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_75 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h4b == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_75 <= 1'h0;
      end else begin
        way1Age_75 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_76 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h4c == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_76 <= 1'h0;
      end else begin
        way1Age_76 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_77 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h4d == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_77 <= 1'h0;
      end else begin
        way1Age_77 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_78 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h4e == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_78 <= 1'h0;
      end else begin
        way1Age_78 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_79 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h4f == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_79 <= 1'h0;
      end else begin
        way1Age_79 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_80 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h50 == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_80 <= 1'h0;
      end else begin
        way1Age_80 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_81 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h51 == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_81 <= 1'h0;
      end else begin
        way1Age_81 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_82 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h52 == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_82 <= 1'h0;
      end else begin
        way1Age_82 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_83 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h53 == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_83 <= 1'h0;
      end else begin
        way1Age_83 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_84 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h54 == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_84 <= 1'h0;
      end else begin
        way1Age_84 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_85 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h55 == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_85 <= 1'h0;
      end else begin
        way1Age_85 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_86 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h56 == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_86 <= 1'h0;
      end else begin
        way1Age_86 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_87 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h57 == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_87 <= 1'h0;
      end else begin
        way1Age_87 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_88 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h58 == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_88 <= 1'h0;
      end else begin
        way1Age_88 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_89 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h59 == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_89 <= 1'h0;
      end else begin
        way1Age_89 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_90 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h5a == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_90 <= 1'h0;
      end else begin
        way1Age_90 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_91 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h5b == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_91 <= 1'h0;
      end else begin
        way1Age_91 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_92 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h5c == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_92 <= 1'h0;
      end else begin
        way1Age_92 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_93 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h5d == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_93 <= 1'h0;
      end else begin
        way1Age_93 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_94 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h5e == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_94 <= 1'h0;
      end else begin
        way1Age_94 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_95 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h5f == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_95 <= 1'h0;
      end else begin
        way1Age_95 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_96 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h60 == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_96 <= 1'h0;
      end else begin
        way1Age_96 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_97 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h61 == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_97 <= 1'h0;
      end else begin
        way1Age_97 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_98 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h62 == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_98 <= 1'h0;
      end else begin
        way1Age_98 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_99 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h63 == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_99 <= 1'h0;
      end else begin
        way1Age_99 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_100 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h64 == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_100 <= 1'h0;
      end else begin
        way1Age_100 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_101 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h65 == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_101 <= 1'h0;
      end else begin
        way1Age_101 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_102 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h66 == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_102 <= 1'h0;
      end else begin
        way1Age_102 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_103 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h67 == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_103 <= 1'h0;
      end else begin
        way1Age_103 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_104 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h68 == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_104 <= 1'h0;
      end else begin
        way1Age_104 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_105 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h69 == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_105 <= 1'h0;
      end else begin
        way1Age_105 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_106 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h6a == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_106 <= 1'h0;
      end else begin
        way1Age_106 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_107 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h6b == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_107 <= 1'h0;
      end else begin
        way1Age_107 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_108 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h6c == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_108 <= 1'h0;
      end else begin
        way1Age_108 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_109 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h6d == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_109 <= 1'h0;
      end else begin
        way1Age_109 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_110 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h6e == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_110 <= 1'h0;
      end else begin
        way1Age_110 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_111 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h6f == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_111 <= 1'h0;
      end else begin
        way1Age_111 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_112 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h70 == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_112 <= 1'h0;
      end else begin
        way1Age_112 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_113 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h71 == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_113 <= 1'h0;
      end else begin
        way1Age_113 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_114 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h72 == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_114 <= 1'h0;
      end else begin
        way1Age_114 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_115 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h73 == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_115 <= 1'h0;
      end else begin
        way1Age_115 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_116 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h74 == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_116 <= 1'h0;
      end else begin
        way1Age_116 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_117 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h75 == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_117 <= 1'h0;
      end else begin
        way1Age_117 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_118 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h76 == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_118 <= 1'h0;
      end else begin
        way1Age_118 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_119 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h77 == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_119 <= 1'h0;
      end else begin
        way1Age_119 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_120 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h78 == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_120 <= 1'h0;
      end else begin
        way1Age_120 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_121 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h79 == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_121 <= 1'h0;
      end else begin
        way1Age_121 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_122 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h7a == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_122 <= 1'h0;
      end else begin
        way1Age_122 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_123 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h7b == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_123 <= 1'h0;
      end else begin
        way1Age_123 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_124 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h7c == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_124 <= 1'h0;
      end else begin
        way1Age_124 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_125 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h7d == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_125 <= 1'h0;
      end else begin
        way1Age_125 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_126 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h7e == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_126 <= 1'h0;
      end else begin
        way1Age_126 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 35:24]
      way1Age_127 <= 1'h0; // @[ICache.scala 35:24]
    end else if (7'h7f == reqIndex) begin // @[ICache.scala 114:21]
      if (ageWay0En) begin // @[ICache.scala 112:25]
        way1Age_127 <= 1'h0;
      end else begin
        way1Age_127 <= 1'h1;
      end
    end
    if (reset) begin // @[ICache.scala 38:22]
      state <= 2'h0; // @[ICache.scala 38:22]
    end else if (2'h0 == state) begin // @[ICache.scala 63:17]
      if (io_imem_inst_valid) begin // @[ICache.scala 65:27]
        state <= 2'h1; // @[ICache.scala 66:15]
      end
    end else if (2'h1 == state) begin // @[ICache.scala 63:17]
      if (cacheHitEn) begin // @[ICache.scala 71:24]
        state <= 2'h0; // @[ICache.scala 72:15]
      end else begin
        state <= 2'h2; // @[ICache.scala 74:15]
      end
    end else if (2'h2 == state) begin // @[ICache.scala 63:17]
      state <= _GEN_514;
    end else begin
      state <= _GEN_515;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {4{`RANDOM}};
  cacheWData = _RAND_0[127:0];
  _RAND_1 = {1{`RANDOM}};
  way0V_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  way0V_1 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  way0V_2 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  way0V_3 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  way0V_4 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  way0V_5 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  way0V_6 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  way0V_7 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  way0V_8 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  way0V_9 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  way0V_10 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  way0V_11 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  way0V_12 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  way0V_13 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  way0V_14 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  way0V_15 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  way0V_16 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  way0V_17 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  way0V_18 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  way0V_19 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  way0V_20 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  way0V_21 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  way0V_22 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  way0V_23 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  way0V_24 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  way0V_25 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  way0V_26 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  way0V_27 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  way0V_28 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  way0V_29 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  way0V_30 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  way0V_31 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  way0V_32 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  way0V_33 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  way0V_34 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  way0V_35 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  way0V_36 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  way0V_37 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  way0V_38 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  way0V_39 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  way0V_40 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  way0V_41 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  way0V_42 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  way0V_43 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  way0V_44 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  way0V_45 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  way0V_46 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  way0V_47 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  way0V_48 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  way0V_49 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  way0V_50 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  way0V_51 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  way0V_52 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  way0V_53 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  way0V_54 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  way0V_55 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  way0V_56 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  way0V_57 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  way0V_58 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  way0V_59 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  way0V_60 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  way0V_61 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  way0V_62 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  way0V_63 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  way0V_64 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  way0V_65 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  way0V_66 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  way0V_67 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  way0V_68 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  way0V_69 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  way0V_70 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  way0V_71 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  way0V_72 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  way0V_73 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  way0V_74 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  way0V_75 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  way0V_76 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  way0V_77 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  way0V_78 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  way0V_79 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  way0V_80 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  way0V_81 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  way0V_82 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  way0V_83 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  way0V_84 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  way0V_85 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  way0V_86 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  way0V_87 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  way0V_88 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  way0V_89 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  way0V_90 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  way0V_91 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  way0V_92 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  way0V_93 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  way0V_94 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  way0V_95 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  way0V_96 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  way0V_97 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  way0V_98 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  way0V_99 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  way0V_100 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  way0V_101 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  way0V_102 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  way0V_103 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  way0V_104 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  way0V_105 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  way0V_106 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  way0V_107 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  way0V_108 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  way0V_109 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  way0V_110 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  way0V_111 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  way0V_112 = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  way0V_113 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  way0V_114 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  way0V_115 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  way0V_116 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  way0V_117 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  way0V_118 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  way0V_119 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  way0V_120 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  way0V_121 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  way0V_122 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  way0V_123 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  way0V_124 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  way0V_125 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  way0V_126 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  way0V_127 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  way0Tag_0 = _RAND_129[20:0];
  _RAND_130 = {1{`RANDOM}};
  way0Tag_1 = _RAND_130[20:0];
  _RAND_131 = {1{`RANDOM}};
  way0Tag_2 = _RAND_131[20:0];
  _RAND_132 = {1{`RANDOM}};
  way0Tag_3 = _RAND_132[20:0];
  _RAND_133 = {1{`RANDOM}};
  way0Tag_4 = _RAND_133[20:0];
  _RAND_134 = {1{`RANDOM}};
  way0Tag_5 = _RAND_134[20:0];
  _RAND_135 = {1{`RANDOM}};
  way0Tag_6 = _RAND_135[20:0];
  _RAND_136 = {1{`RANDOM}};
  way0Tag_7 = _RAND_136[20:0];
  _RAND_137 = {1{`RANDOM}};
  way0Tag_8 = _RAND_137[20:0];
  _RAND_138 = {1{`RANDOM}};
  way0Tag_9 = _RAND_138[20:0];
  _RAND_139 = {1{`RANDOM}};
  way0Tag_10 = _RAND_139[20:0];
  _RAND_140 = {1{`RANDOM}};
  way0Tag_11 = _RAND_140[20:0];
  _RAND_141 = {1{`RANDOM}};
  way0Tag_12 = _RAND_141[20:0];
  _RAND_142 = {1{`RANDOM}};
  way0Tag_13 = _RAND_142[20:0];
  _RAND_143 = {1{`RANDOM}};
  way0Tag_14 = _RAND_143[20:0];
  _RAND_144 = {1{`RANDOM}};
  way0Tag_15 = _RAND_144[20:0];
  _RAND_145 = {1{`RANDOM}};
  way0Tag_16 = _RAND_145[20:0];
  _RAND_146 = {1{`RANDOM}};
  way0Tag_17 = _RAND_146[20:0];
  _RAND_147 = {1{`RANDOM}};
  way0Tag_18 = _RAND_147[20:0];
  _RAND_148 = {1{`RANDOM}};
  way0Tag_19 = _RAND_148[20:0];
  _RAND_149 = {1{`RANDOM}};
  way0Tag_20 = _RAND_149[20:0];
  _RAND_150 = {1{`RANDOM}};
  way0Tag_21 = _RAND_150[20:0];
  _RAND_151 = {1{`RANDOM}};
  way0Tag_22 = _RAND_151[20:0];
  _RAND_152 = {1{`RANDOM}};
  way0Tag_23 = _RAND_152[20:0];
  _RAND_153 = {1{`RANDOM}};
  way0Tag_24 = _RAND_153[20:0];
  _RAND_154 = {1{`RANDOM}};
  way0Tag_25 = _RAND_154[20:0];
  _RAND_155 = {1{`RANDOM}};
  way0Tag_26 = _RAND_155[20:0];
  _RAND_156 = {1{`RANDOM}};
  way0Tag_27 = _RAND_156[20:0];
  _RAND_157 = {1{`RANDOM}};
  way0Tag_28 = _RAND_157[20:0];
  _RAND_158 = {1{`RANDOM}};
  way0Tag_29 = _RAND_158[20:0];
  _RAND_159 = {1{`RANDOM}};
  way0Tag_30 = _RAND_159[20:0];
  _RAND_160 = {1{`RANDOM}};
  way0Tag_31 = _RAND_160[20:0];
  _RAND_161 = {1{`RANDOM}};
  way0Tag_32 = _RAND_161[20:0];
  _RAND_162 = {1{`RANDOM}};
  way0Tag_33 = _RAND_162[20:0];
  _RAND_163 = {1{`RANDOM}};
  way0Tag_34 = _RAND_163[20:0];
  _RAND_164 = {1{`RANDOM}};
  way0Tag_35 = _RAND_164[20:0];
  _RAND_165 = {1{`RANDOM}};
  way0Tag_36 = _RAND_165[20:0];
  _RAND_166 = {1{`RANDOM}};
  way0Tag_37 = _RAND_166[20:0];
  _RAND_167 = {1{`RANDOM}};
  way0Tag_38 = _RAND_167[20:0];
  _RAND_168 = {1{`RANDOM}};
  way0Tag_39 = _RAND_168[20:0];
  _RAND_169 = {1{`RANDOM}};
  way0Tag_40 = _RAND_169[20:0];
  _RAND_170 = {1{`RANDOM}};
  way0Tag_41 = _RAND_170[20:0];
  _RAND_171 = {1{`RANDOM}};
  way0Tag_42 = _RAND_171[20:0];
  _RAND_172 = {1{`RANDOM}};
  way0Tag_43 = _RAND_172[20:0];
  _RAND_173 = {1{`RANDOM}};
  way0Tag_44 = _RAND_173[20:0];
  _RAND_174 = {1{`RANDOM}};
  way0Tag_45 = _RAND_174[20:0];
  _RAND_175 = {1{`RANDOM}};
  way0Tag_46 = _RAND_175[20:0];
  _RAND_176 = {1{`RANDOM}};
  way0Tag_47 = _RAND_176[20:0];
  _RAND_177 = {1{`RANDOM}};
  way0Tag_48 = _RAND_177[20:0];
  _RAND_178 = {1{`RANDOM}};
  way0Tag_49 = _RAND_178[20:0];
  _RAND_179 = {1{`RANDOM}};
  way0Tag_50 = _RAND_179[20:0];
  _RAND_180 = {1{`RANDOM}};
  way0Tag_51 = _RAND_180[20:0];
  _RAND_181 = {1{`RANDOM}};
  way0Tag_52 = _RAND_181[20:0];
  _RAND_182 = {1{`RANDOM}};
  way0Tag_53 = _RAND_182[20:0];
  _RAND_183 = {1{`RANDOM}};
  way0Tag_54 = _RAND_183[20:0];
  _RAND_184 = {1{`RANDOM}};
  way0Tag_55 = _RAND_184[20:0];
  _RAND_185 = {1{`RANDOM}};
  way0Tag_56 = _RAND_185[20:0];
  _RAND_186 = {1{`RANDOM}};
  way0Tag_57 = _RAND_186[20:0];
  _RAND_187 = {1{`RANDOM}};
  way0Tag_58 = _RAND_187[20:0];
  _RAND_188 = {1{`RANDOM}};
  way0Tag_59 = _RAND_188[20:0];
  _RAND_189 = {1{`RANDOM}};
  way0Tag_60 = _RAND_189[20:0];
  _RAND_190 = {1{`RANDOM}};
  way0Tag_61 = _RAND_190[20:0];
  _RAND_191 = {1{`RANDOM}};
  way0Tag_62 = _RAND_191[20:0];
  _RAND_192 = {1{`RANDOM}};
  way0Tag_63 = _RAND_192[20:0];
  _RAND_193 = {1{`RANDOM}};
  way0Tag_64 = _RAND_193[20:0];
  _RAND_194 = {1{`RANDOM}};
  way0Tag_65 = _RAND_194[20:0];
  _RAND_195 = {1{`RANDOM}};
  way0Tag_66 = _RAND_195[20:0];
  _RAND_196 = {1{`RANDOM}};
  way0Tag_67 = _RAND_196[20:0];
  _RAND_197 = {1{`RANDOM}};
  way0Tag_68 = _RAND_197[20:0];
  _RAND_198 = {1{`RANDOM}};
  way0Tag_69 = _RAND_198[20:0];
  _RAND_199 = {1{`RANDOM}};
  way0Tag_70 = _RAND_199[20:0];
  _RAND_200 = {1{`RANDOM}};
  way0Tag_71 = _RAND_200[20:0];
  _RAND_201 = {1{`RANDOM}};
  way0Tag_72 = _RAND_201[20:0];
  _RAND_202 = {1{`RANDOM}};
  way0Tag_73 = _RAND_202[20:0];
  _RAND_203 = {1{`RANDOM}};
  way0Tag_74 = _RAND_203[20:0];
  _RAND_204 = {1{`RANDOM}};
  way0Tag_75 = _RAND_204[20:0];
  _RAND_205 = {1{`RANDOM}};
  way0Tag_76 = _RAND_205[20:0];
  _RAND_206 = {1{`RANDOM}};
  way0Tag_77 = _RAND_206[20:0];
  _RAND_207 = {1{`RANDOM}};
  way0Tag_78 = _RAND_207[20:0];
  _RAND_208 = {1{`RANDOM}};
  way0Tag_79 = _RAND_208[20:0];
  _RAND_209 = {1{`RANDOM}};
  way0Tag_80 = _RAND_209[20:0];
  _RAND_210 = {1{`RANDOM}};
  way0Tag_81 = _RAND_210[20:0];
  _RAND_211 = {1{`RANDOM}};
  way0Tag_82 = _RAND_211[20:0];
  _RAND_212 = {1{`RANDOM}};
  way0Tag_83 = _RAND_212[20:0];
  _RAND_213 = {1{`RANDOM}};
  way0Tag_84 = _RAND_213[20:0];
  _RAND_214 = {1{`RANDOM}};
  way0Tag_85 = _RAND_214[20:0];
  _RAND_215 = {1{`RANDOM}};
  way0Tag_86 = _RAND_215[20:0];
  _RAND_216 = {1{`RANDOM}};
  way0Tag_87 = _RAND_216[20:0];
  _RAND_217 = {1{`RANDOM}};
  way0Tag_88 = _RAND_217[20:0];
  _RAND_218 = {1{`RANDOM}};
  way0Tag_89 = _RAND_218[20:0];
  _RAND_219 = {1{`RANDOM}};
  way0Tag_90 = _RAND_219[20:0];
  _RAND_220 = {1{`RANDOM}};
  way0Tag_91 = _RAND_220[20:0];
  _RAND_221 = {1{`RANDOM}};
  way0Tag_92 = _RAND_221[20:0];
  _RAND_222 = {1{`RANDOM}};
  way0Tag_93 = _RAND_222[20:0];
  _RAND_223 = {1{`RANDOM}};
  way0Tag_94 = _RAND_223[20:0];
  _RAND_224 = {1{`RANDOM}};
  way0Tag_95 = _RAND_224[20:0];
  _RAND_225 = {1{`RANDOM}};
  way0Tag_96 = _RAND_225[20:0];
  _RAND_226 = {1{`RANDOM}};
  way0Tag_97 = _RAND_226[20:0];
  _RAND_227 = {1{`RANDOM}};
  way0Tag_98 = _RAND_227[20:0];
  _RAND_228 = {1{`RANDOM}};
  way0Tag_99 = _RAND_228[20:0];
  _RAND_229 = {1{`RANDOM}};
  way0Tag_100 = _RAND_229[20:0];
  _RAND_230 = {1{`RANDOM}};
  way0Tag_101 = _RAND_230[20:0];
  _RAND_231 = {1{`RANDOM}};
  way0Tag_102 = _RAND_231[20:0];
  _RAND_232 = {1{`RANDOM}};
  way0Tag_103 = _RAND_232[20:0];
  _RAND_233 = {1{`RANDOM}};
  way0Tag_104 = _RAND_233[20:0];
  _RAND_234 = {1{`RANDOM}};
  way0Tag_105 = _RAND_234[20:0];
  _RAND_235 = {1{`RANDOM}};
  way0Tag_106 = _RAND_235[20:0];
  _RAND_236 = {1{`RANDOM}};
  way0Tag_107 = _RAND_236[20:0];
  _RAND_237 = {1{`RANDOM}};
  way0Tag_108 = _RAND_237[20:0];
  _RAND_238 = {1{`RANDOM}};
  way0Tag_109 = _RAND_238[20:0];
  _RAND_239 = {1{`RANDOM}};
  way0Tag_110 = _RAND_239[20:0];
  _RAND_240 = {1{`RANDOM}};
  way0Tag_111 = _RAND_240[20:0];
  _RAND_241 = {1{`RANDOM}};
  way0Tag_112 = _RAND_241[20:0];
  _RAND_242 = {1{`RANDOM}};
  way0Tag_113 = _RAND_242[20:0];
  _RAND_243 = {1{`RANDOM}};
  way0Tag_114 = _RAND_243[20:0];
  _RAND_244 = {1{`RANDOM}};
  way0Tag_115 = _RAND_244[20:0];
  _RAND_245 = {1{`RANDOM}};
  way0Tag_116 = _RAND_245[20:0];
  _RAND_246 = {1{`RANDOM}};
  way0Tag_117 = _RAND_246[20:0];
  _RAND_247 = {1{`RANDOM}};
  way0Tag_118 = _RAND_247[20:0];
  _RAND_248 = {1{`RANDOM}};
  way0Tag_119 = _RAND_248[20:0];
  _RAND_249 = {1{`RANDOM}};
  way0Tag_120 = _RAND_249[20:0];
  _RAND_250 = {1{`RANDOM}};
  way0Tag_121 = _RAND_250[20:0];
  _RAND_251 = {1{`RANDOM}};
  way0Tag_122 = _RAND_251[20:0];
  _RAND_252 = {1{`RANDOM}};
  way0Tag_123 = _RAND_252[20:0];
  _RAND_253 = {1{`RANDOM}};
  way0Tag_124 = _RAND_253[20:0];
  _RAND_254 = {1{`RANDOM}};
  way0Tag_125 = _RAND_254[20:0];
  _RAND_255 = {1{`RANDOM}};
  way0Tag_126 = _RAND_255[20:0];
  _RAND_256 = {1{`RANDOM}};
  way0Tag_127 = _RAND_256[20:0];
  _RAND_257 = {1{`RANDOM}};
  way0Age_0 = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  way0Age_1 = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  way0Age_2 = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  way0Age_3 = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  way0Age_4 = _RAND_261[0:0];
  _RAND_262 = {1{`RANDOM}};
  way0Age_5 = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  way0Age_6 = _RAND_263[0:0];
  _RAND_264 = {1{`RANDOM}};
  way0Age_7 = _RAND_264[0:0];
  _RAND_265 = {1{`RANDOM}};
  way0Age_8 = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  way0Age_9 = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  way0Age_10 = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  way0Age_11 = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  way0Age_12 = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  way0Age_13 = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  way0Age_14 = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  way0Age_15 = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  way0Age_16 = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  way0Age_17 = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  way0Age_18 = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  way0Age_19 = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  way0Age_20 = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  way0Age_21 = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  way0Age_22 = _RAND_279[0:0];
  _RAND_280 = {1{`RANDOM}};
  way0Age_23 = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  way0Age_24 = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  way0Age_25 = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  way0Age_26 = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  way0Age_27 = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  way0Age_28 = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  way0Age_29 = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  way0Age_30 = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  way0Age_31 = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  way0Age_32 = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  way0Age_33 = _RAND_290[0:0];
  _RAND_291 = {1{`RANDOM}};
  way0Age_34 = _RAND_291[0:0];
  _RAND_292 = {1{`RANDOM}};
  way0Age_35 = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  way0Age_36 = _RAND_293[0:0];
  _RAND_294 = {1{`RANDOM}};
  way0Age_37 = _RAND_294[0:0];
  _RAND_295 = {1{`RANDOM}};
  way0Age_38 = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  way0Age_39 = _RAND_296[0:0];
  _RAND_297 = {1{`RANDOM}};
  way0Age_40 = _RAND_297[0:0];
  _RAND_298 = {1{`RANDOM}};
  way0Age_41 = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  way0Age_42 = _RAND_299[0:0];
  _RAND_300 = {1{`RANDOM}};
  way0Age_43 = _RAND_300[0:0];
  _RAND_301 = {1{`RANDOM}};
  way0Age_44 = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  way0Age_45 = _RAND_302[0:0];
  _RAND_303 = {1{`RANDOM}};
  way0Age_46 = _RAND_303[0:0];
  _RAND_304 = {1{`RANDOM}};
  way0Age_47 = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  way0Age_48 = _RAND_305[0:0];
  _RAND_306 = {1{`RANDOM}};
  way0Age_49 = _RAND_306[0:0];
  _RAND_307 = {1{`RANDOM}};
  way0Age_50 = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  way0Age_51 = _RAND_308[0:0];
  _RAND_309 = {1{`RANDOM}};
  way0Age_52 = _RAND_309[0:0];
  _RAND_310 = {1{`RANDOM}};
  way0Age_53 = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  way0Age_54 = _RAND_311[0:0];
  _RAND_312 = {1{`RANDOM}};
  way0Age_55 = _RAND_312[0:0];
  _RAND_313 = {1{`RANDOM}};
  way0Age_56 = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  way0Age_57 = _RAND_314[0:0];
  _RAND_315 = {1{`RANDOM}};
  way0Age_58 = _RAND_315[0:0];
  _RAND_316 = {1{`RANDOM}};
  way0Age_59 = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  way0Age_60 = _RAND_317[0:0];
  _RAND_318 = {1{`RANDOM}};
  way0Age_61 = _RAND_318[0:0];
  _RAND_319 = {1{`RANDOM}};
  way0Age_62 = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  way0Age_63 = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  way0Age_64 = _RAND_321[0:0];
  _RAND_322 = {1{`RANDOM}};
  way0Age_65 = _RAND_322[0:0];
  _RAND_323 = {1{`RANDOM}};
  way0Age_66 = _RAND_323[0:0];
  _RAND_324 = {1{`RANDOM}};
  way0Age_67 = _RAND_324[0:0];
  _RAND_325 = {1{`RANDOM}};
  way0Age_68 = _RAND_325[0:0];
  _RAND_326 = {1{`RANDOM}};
  way0Age_69 = _RAND_326[0:0];
  _RAND_327 = {1{`RANDOM}};
  way0Age_70 = _RAND_327[0:0];
  _RAND_328 = {1{`RANDOM}};
  way0Age_71 = _RAND_328[0:0];
  _RAND_329 = {1{`RANDOM}};
  way0Age_72 = _RAND_329[0:0];
  _RAND_330 = {1{`RANDOM}};
  way0Age_73 = _RAND_330[0:0];
  _RAND_331 = {1{`RANDOM}};
  way0Age_74 = _RAND_331[0:0];
  _RAND_332 = {1{`RANDOM}};
  way0Age_75 = _RAND_332[0:0];
  _RAND_333 = {1{`RANDOM}};
  way0Age_76 = _RAND_333[0:0];
  _RAND_334 = {1{`RANDOM}};
  way0Age_77 = _RAND_334[0:0];
  _RAND_335 = {1{`RANDOM}};
  way0Age_78 = _RAND_335[0:0];
  _RAND_336 = {1{`RANDOM}};
  way0Age_79 = _RAND_336[0:0];
  _RAND_337 = {1{`RANDOM}};
  way0Age_80 = _RAND_337[0:0];
  _RAND_338 = {1{`RANDOM}};
  way0Age_81 = _RAND_338[0:0];
  _RAND_339 = {1{`RANDOM}};
  way0Age_82 = _RAND_339[0:0];
  _RAND_340 = {1{`RANDOM}};
  way0Age_83 = _RAND_340[0:0];
  _RAND_341 = {1{`RANDOM}};
  way0Age_84 = _RAND_341[0:0];
  _RAND_342 = {1{`RANDOM}};
  way0Age_85 = _RAND_342[0:0];
  _RAND_343 = {1{`RANDOM}};
  way0Age_86 = _RAND_343[0:0];
  _RAND_344 = {1{`RANDOM}};
  way0Age_87 = _RAND_344[0:0];
  _RAND_345 = {1{`RANDOM}};
  way0Age_88 = _RAND_345[0:0];
  _RAND_346 = {1{`RANDOM}};
  way0Age_89 = _RAND_346[0:0];
  _RAND_347 = {1{`RANDOM}};
  way0Age_90 = _RAND_347[0:0];
  _RAND_348 = {1{`RANDOM}};
  way0Age_91 = _RAND_348[0:0];
  _RAND_349 = {1{`RANDOM}};
  way0Age_92 = _RAND_349[0:0];
  _RAND_350 = {1{`RANDOM}};
  way0Age_93 = _RAND_350[0:0];
  _RAND_351 = {1{`RANDOM}};
  way0Age_94 = _RAND_351[0:0];
  _RAND_352 = {1{`RANDOM}};
  way0Age_95 = _RAND_352[0:0];
  _RAND_353 = {1{`RANDOM}};
  way0Age_96 = _RAND_353[0:0];
  _RAND_354 = {1{`RANDOM}};
  way0Age_97 = _RAND_354[0:0];
  _RAND_355 = {1{`RANDOM}};
  way0Age_98 = _RAND_355[0:0];
  _RAND_356 = {1{`RANDOM}};
  way0Age_99 = _RAND_356[0:0];
  _RAND_357 = {1{`RANDOM}};
  way0Age_100 = _RAND_357[0:0];
  _RAND_358 = {1{`RANDOM}};
  way0Age_101 = _RAND_358[0:0];
  _RAND_359 = {1{`RANDOM}};
  way0Age_102 = _RAND_359[0:0];
  _RAND_360 = {1{`RANDOM}};
  way0Age_103 = _RAND_360[0:0];
  _RAND_361 = {1{`RANDOM}};
  way0Age_104 = _RAND_361[0:0];
  _RAND_362 = {1{`RANDOM}};
  way0Age_105 = _RAND_362[0:0];
  _RAND_363 = {1{`RANDOM}};
  way0Age_106 = _RAND_363[0:0];
  _RAND_364 = {1{`RANDOM}};
  way0Age_107 = _RAND_364[0:0];
  _RAND_365 = {1{`RANDOM}};
  way0Age_108 = _RAND_365[0:0];
  _RAND_366 = {1{`RANDOM}};
  way0Age_109 = _RAND_366[0:0];
  _RAND_367 = {1{`RANDOM}};
  way0Age_110 = _RAND_367[0:0];
  _RAND_368 = {1{`RANDOM}};
  way0Age_111 = _RAND_368[0:0];
  _RAND_369 = {1{`RANDOM}};
  way0Age_112 = _RAND_369[0:0];
  _RAND_370 = {1{`RANDOM}};
  way0Age_113 = _RAND_370[0:0];
  _RAND_371 = {1{`RANDOM}};
  way0Age_114 = _RAND_371[0:0];
  _RAND_372 = {1{`RANDOM}};
  way0Age_115 = _RAND_372[0:0];
  _RAND_373 = {1{`RANDOM}};
  way0Age_116 = _RAND_373[0:0];
  _RAND_374 = {1{`RANDOM}};
  way0Age_117 = _RAND_374[0:0];
  _RAND_375 = {1{`RANDOM}};
  way0Age_118 = _RAND_375[0:0];
  _RAND_376 = {1{`RANDOM}};
  way0Age_119 = _RAND_376[0:0];
  _RAND_377 = {1{`RANDOM}};
  way0Age_120 = _RAND_377[0:0];
  _RAND_378 = {1{`RANDOM}};
  way0Age_121 = _RAND_378[0:0];
  _RAND_379 = {1{`RANDOM}};
  way0Age_122 = _RAND_379[0:0];
  _RAND_380 = {1{`RANDOM}};
  way0Age_123 = _RAND_380[0:0];
  _RAND_381 = {1{`RANDOM}};
  way0Age_124 = _RAND_381[0:0];
  _RAND_382 = {1{`RANDOM}};
  way0Age_125 = _RAND_382[0:0];
  _RAND_383 = {1{`RANDOM}};
  way0Age_126 = _RAND_383[0:0];
  _RAND_384 = {1{`RANDOM}};
  way0Age_127 = _RAND_384[0:0];
  _RAND_385 = {1{`RANDOM}};
  way1V_0 = _RAND_385[0:0];
  _RAND_386 = {1{`RANDOM}};
  way1V_1 = _RAND_386[0:0];
  _RAND_387 = {1{`RANDOM}};
  way1V_2 = _RAND_387[0:0];
  _RAND_388 = {1{`RANDOM}};
  way1V_3 = _RAND_388[0:0];
  _RAND_389 = {1{`RANDOM}};
  way1V_4 = _RAND_389[0:0];
  _RAND_390 = {1{`RANDOM}};
  way1V_5 = _RAND_390[0:0];
  _RAND_391 = {1{`RANDOM}};
  way1V_6 = _RAND_391[0:0];
  _RAND_392 = {1{`RANDOM}};
  way1V_7 = _RAND_392[0:0];
  _RAND_393 = {1{`RANDOM}};
  way1V_8 = _RAND_393[0:0];
  _RAND_394 = {1{`RANDOM}};
  way1V_9 = _RAND_394[0:0];
  _RAND_395 = {1{`RANDOM}};
  way1V_10 = _RAND_395[0:0];
  _RAND_396 = {1{`RANDOM}};
  way1V_11 = _RAND_396[0:0];
  _RAND_397 = {1{`RANDOM}};
  way1V_12 = _RAND_397[0:0];
  _RAND_398 = {1{`RANDOM}};
  way1V_13 = _RAND_398[0:0];
  _RAND_399 = {1{`RANDOM}};
  way1V_14 = _RAND_399[0:0];
  _RAND_400 = {1{`RANDOM}};
  way1V_15 = _RAND_400[0:0];
  _RAND_401 = {1{`RANDOM}};
  way1V_16 = _RAND_401[0:0];
  _RAND_402 = {1{`RANDOM}};
  way1V_17 = _RAND_402[0:0];
  _RAND_403 = {1{`RANDOM}};
  way1V_18 = _RAND_403[0:0];
  _RAND_404 = {1{`RANDOM}};
  way1V_19 = _RAND_404[0:0];
  _RAND_405 = {1{`RANDOM}};
  way1V_20 = _RAND_405[0:0];
  _RAND_406 = {1{`RANDOM}};
  way1V_21 = _RAND_406[0:0];
  _RAND_407 = {1{`RANDOM}};
  way1V_22 = _RAND_407[0:0];
  _RAND_408 = {1{`RANDOM}};
  way1V_23 = _RAND_408[0:0];
  _RAND_409 = {1{`RANDOM}};
  way1V_24 = _RAND_409[0:0];
  _RAND_410 = {1{`RANDOM}};
  way1V_25 = _RAND_410[0:0];
  _RAND_411 = {1{`RANDOM}};
  way1V_26 = _RAND_411[0:0];
  _RAND_412 = {1{`RANDOM}};
  way1V_27 = _RAND_412[0:0];
  _RAND_413 = {1{`RANDOM}};
  way1V_28 = _RAND_413[0:0];
  _RAND_414 = {1{`RANDOM}};
  way1V_29 = _RAND_414[0:0];
  _RAND_415 = {1{`RANDOM}};
  way1V_30 = _RAND_415[0:0];
  _RAND_416 = {1{`RANDOM}};
  way1V_31 = _RAND_416[0:0];
  _RAND_417 = {1{`RANDOM}};
  way1V_32 = _RAND_417[0:0];
  _RAND_418 = {1{`RANDOM}};
  way1V_33 = _RAND_418[0:0];
  _RAND_419 = {1{`RANDOM}};
  way1V_34 = _RAND_419[0:0];
  _RAND_420 = {1{`RANDOM}};
  way1V_35 = _RAND_420[0:0];
  _RAND_421 = {1{`RANDOM}};
  way1V_36 = _RAND_421[0:0];
  _RAND_422 = {1{`RANDOM}};
  way1V_37 = _RAND_422[0:0];
  _RAND_423 = {1{`RANDOM}};
  way1V_38 = _RAND_423[0:0];
  _RAND_424 = {1{`RANDOM}};
  way1V_39 = _RAND_424[0:0];
  _RAND_425 = {1{`RANDOM}};
  way1V_40 = _RAND_425[0:0];
  _RAND_426 = {1{`RANDOM}};
  way1V_41 = _RAND_426[0:0];
  _RAND_427 = {1{`RANDOM}};
  way1V_42 = _RAND_427[0:0];
  _RAND_428 = {1{`RANDOM}};
  way1V_43 = _RAND_428[0:0];
  _RAND_429 = {1{`RANDOM}};
  way1V_44 = _RAND_429[0:0];
  _RAND_430 = {1{`RANDOM}};
  way1V_45 = _RAND_430[0:0];
  _RAND_431 = {1{`RANDOM}};
  way1V_46 = _RAND_431[0:0];
  _RAND_432 = {1{`RANDOM}};
  way1V_47 = _RAND_432[0:0];
  _RAND_433 = {1{`RANDOM}};
  way1V_48 = _RAND_433[0:0];
  _RAND_434 = {1{`RANDOM}};
  way1V_49 = _RAND_434[0:0];
  _RAND_435 = {1{`RANDOM}};
  way1V_50 = _RAND_435[0:0];
  _RAND_436 = {1{`RANDOM}};
  way1V_51 = _RAND_436[0:0];
  _RAND_437 = {1{`RANDOM}};
  way1V_52 = _RAND_437[0:0];
  _RAND_438 = {1{`RANDOM}};
  way1V_53 = _RAND_438[0:0];
  _RAND_439 = {1{`RANDOM}};
  way1V_54 = _RAND_439[0:0];
  _RAND_440 = {1{`RANDOM}};
  way1V_55 = _RAND_440[0:0];
  _RAND_441 = {1{`RANDOM}};
  way1V_56 = _RAND_441[0:0];
  _RAND_442 = {1{`RANDOM}};
  way1V_57 = _RAND_442[0:0];
  _RAND_443 = {1{`RANDOM}};
  way1V_58 = _RAND_443[0:0];
  _RAND_444 = {1{`RANDOM}};
  way1V_59 = _RAND_444[0:0];
  _RAND_445 = {1{`RANDOM}};
  way1V_60 = _RAND_445[0:0];
  _RAND_446 = {1{`RANDOM}};
  way1V_61 = _RAND_446[0:0];
  _RAND_447 = {1{`RANDOM}};
  way1V_62 = _RAND_447[0:0];
  _RAND_448 = {1{`RANDOM}};
  way1V_63 = _RAND_448[0:0];
  _RAND_449 = {1{`RANDOM}};
  way1V_64 = _RAND_449[0:0];
  _RAND_450 = {1{`RANDOM}};
  way1V_65 = _RAND_450[0:0];
  _RAND_451 = {1{`RANDOM}};
  way1V_66 = _RAND_451[0:0];
  _RAND_452 = {1{`RANDOM}};
  way1V_67 = _RAND_452[0:0];
  _RAND_453 = {1{`RANDOM}};
  way1V_68 = _RAND_453[0:0];
  _RAND_454 = {1{`RANDOM}};
  way1V_69 = _RAND_454[0:0];
  _RAND_455 = {1{`RANDOM}};
  way1V_70 = _RAND_455[0:0];
  _RAND_456 = {1{`RANDOM}};
  way1V_71 = _RAND_456[0:0];
  _RAND_457 = {1{`RANDOM}};
  way1V_72 = _RAND_457[0:0];
  _RAND_458 = {1{`RANDOM}};
  way1V_73 = _RAND_458[0:0];
  _RAND_459 = {1{`RANDOM}};
  way1V_74 = _RAND_459[0:0];
  _RAND_460 = {1{`RANDOM}};
  way1V_75 = _RAND_460[0:0];
  _RAND_461 = {1{`RANDOM}};
  way1V_76 = _RAND_461[0:0];
  _RAND_462 = {1{`RANDOM}};
  way1V_77 = _RAND_462[0:0];
  _RAND_463 = {1{`RANDOM}};
  way1V_78 = _RAND_463[0:0];
  _RAND_464 = {1{`RANDOM}};
  way1V_79 = _RAND_464[0:0];
  _RAND_465 = {1{`RANDOM}};
  way1V_80 = _RAND_465[0:0];
  _RAND_466 = {1{`RANDOM}};
  way1V_81 = _RAND_466[0:0];
  _RAND_467 = {1{`RANDOM}};
  way1V_82 = _RAND_467[0:0];
  _RAND_468 = {1{`RANDOM}};
  way1V_83 = _RAND_468[0:0];
  _RAND_469 = {1{`RANDOM}};
  way1V_84 = _RAND_469[0:0];
  _RAND_470 = {1{`RANDOM}};
  way1V_85 = _RAND_470[0:0];
  _RAND_471 = {1{`RANDOM}};
  way1V_86 = _RAND_471[0:0];
  _RAND_472 = {1{`RANDOM}};
  way1V_87 = _RAND_472[0:0];
  _RAND_473 = {1{`RANDOM}};
  way1V_88 = _RAND_473[0:0];
  _RAND_474 = {1{`RANDOM}};
  way1V_89 = _RAND_474[0:0];
  _RAND_475 = {1{`RANDOM}};
  way1V_90 = _RAND_475[0:0];
  _RAND_476 = {1{`RANDOM}};
  way1V_91 = _RAND_476[0:0];
  _RAND_477 = {1{`RANDOM}};
  way1V_92 = _RAND_477[0:0];
  _RAND_478 = {1{`RANDOM}};
  way1V_93 = _RAND_478[0:0];
  _RAND_479 = {1{`RANDOM}};
  way1V_94 = _RAND_479[0:0];
  _RAND_480 = {1{`RANDOM}};
  way1V_95 = _RAND_480[0:0];
  _RAND_481 = {1{`RANDOM}};
  way1V_96 = _RAND_481[0:0];
  _RAND_482 = {1{`RANDOM}};
  way1V_97 = _RAND_482[0:0];
  _RAND_483 = {1{`RANDOM}};
  way1V_98 = _RAND_483[0:0];
  _RAND_484 = {1{`RANDOM}};
  way1V_99 = _RAND_484[0:0];
  _RAND_485 = {1{`RANDOM}};
  way1V_100 = _RAND_485[0:0];
  _RAND_486 = {1{`RANDOM}};
  way1V_101 = _RAND_486[0:0];
  _RAND_487 = {1{`RANDOM}};
  way1V_102 = _RAND_487[0:0];
  _RAND_488 = {1{`RANDOM}};
  way1V_103 = _RAND_488[0:0];
  _RAND_489 = {1{`RANDOM}};
  way1V_104 = _RAND_489[0:0];
  _RAND_490 = {1{`RANDOM}};
  way1V_105 = _RAND_490[0:0];
  _RAND_491 = {1{`RANDOM}};
  way1V_106 = _RAND_491[0:0];
  _RAND_492 = {1{`RANDOM}};
  way1V_107 = _RAND_492[0:0];
  _RAND_493 = {1{`RANDOM}};
  way1V_108 = _RAND_493[0:0];
  _RAND_494 = {1{`RANDOM}};
  way1V_109 = _RAND_494[0:0];
  _RAND_495 = {1{`RANDOM}};
  way1V_110 = _RAND_495[0:0];
  _RAND_496 = {1{`RANDOM}};
  way1V_111 = _RAND_496[0:0];
  _RAND_497 = {1{`RANDOM}};
  way1V_112 = _RAND_497[0:0];
  _RAND_498 = {1{`RANDOM}};
  way1V_113 = _RAND_498[0:0];
  _RAND_499 = {1{`RANDOM}};
  way1V_114 = _RAND_499[0:0];
  _RAND_500 = {1{`RANDOM}};
  way1V_115 = _RAND_500[0:0];
  _RAND_501 = {1{`RANDOM}};
  way1V_116 = _RAND_501[0:0];
  _RAND_502 = {1{`RANDOM}};
  way1V_117 = _RAND_502[0:0];
  _RAND_503 = {1{`RANDOM}};
  way1V_118 = _RAND_503[0:0];
  _RAND_504 = {1{`RANDOM}};
  way1V_119 = _RAND_504[0:0];
  _RAND_505 = {1{`RANDOM}};
  way1V_120 = _RAND_505[0:0];
  _RAND_506 = {1{`RANDOM}};
  way1V_121 = _RAND_506[0:0];
  _RAND_507 = {1{`RANDOM}};
  way1V_122 = _RAND_507[0:0];
  _RAND_508 = {1{`RANDOM}};
  way1V_123 = _RAND_508[0:0];
  _RAND_509 = {1{`RANDOM}};
  way1V_124 = _RAND_509[0:0];
  _RAND_510 = {1{`RANDOM}};
  way1V_125 = _RAND_510[0:0];
  _RAND_511 = {1{`RANDOM}};
  way1V_126 = _RAND_511[0:0];
  _RAND_512 = {1{`RANDOM}};
  way1V_127 = _RAND_512[0:0];
  _RAND_513 = {1{`RANDOM}};
  way1Tag_0 = _RAND_513[20:0];
  _RAND_514 = {1{`RANDOM}};
  way1Tag_1 = _RAND_514[20:0];
  _RAND_515 = {1{`RANDOM}};
  way1Tag_2 = _RAND_515[20:0];
  _RAND_516 = {1{`RANDOM}};
  way1Tag_3 = _RAND_516[20:0];
  _RAND_517 = {1{`RANDOM}};
  way1Tag_4 = _RAND_517[20:0];
  _RAND_518 = {1{`RANDOM}};
  way1Tag_5 = _RAND_518[20:0];
  _RAND_519 = {1{`RANDOM}};
  way1Tag_6 = _RAND_519[20:0];
  _RAND_520 = {1{`RANDOM}};
  way1Tag_7 = _RAND_520[20:0];
  _RAND_521 = {1{`RANDOM}};
  way1Tag_8 = _RAND_521[20:0];
  _RAND_522 = {1{`RANDOM}};
  way1Tag_9 = _RAND_522[20:0];
  _RAND_523 = {1{`RANDOM}};
  way1Tag_10 = _RAND_523[20:0];
  _RAND_524 = {1{`RANDOM}};
  way1Tag_11 = _RAND_524[20:0];
  _RAND_525 = {1{`RANDOM}};
  way1Tag_12 = _RAND_525[20:0];
  _RAND_526 = {1{`RANDOM}};
  way1Tag_13 = _RAND_526[20:0];
  _RAND_527 = {1{`RANDOM}};
  way1Tag_14 = _RAND_527[20:0];
  _RAND_528 = {1{`RANDOM}};
  way1Tag_15 = _RAND_528[20:0];
  _RAND_529 = {1{`RANDOM}};
  way1Tag_16 = _RAND_529[20:0];
  _RAND_530 = {1{`RANDOM}};
  way1Tag_17 = _RAND_530[20:0];
  _RAND_531 = {1{`RANDOM}};
  way1Tag_18 = _RAND_531[20:0];
  _RAND_532 = {1{`RANDOM}};
  way1Tag_19 = _RAND_532[20:0];
  _RAND_533 = {1{`RANDOM}};
  way1Tag_20 = _RAND_533[20:0];
  _RAND_534 = {1{`RANDOM}};
  way1Tag_21 = _RAND_534[20:0];
  _RAND_535 = {1{`RANDOM}};
  way1Tag_22 = _RAND_535[20:0];
  _RAND_536 = {1{`RANDOM}};
  way1Tag_23 = _RAND_536[20:0];
  _RAND_537 = {1{`RANDOM}};
  way1Tag_24 = _RAND_537[20:0];
  _RAND_538 = {1{`RANDOM}};
  way1Tag_25 = _RAND_538[20:0];
  _RAND_539 = {1{`RANDOM}};
  way1Tag_26 = _RAND_539[20:0];
  _RAND_540 = {1{`RANDOM}};
  way1Tag_27 = _RAND_540[20:0];
  _RAND_541 = {1{`RANDOM}};
  way1Tag_28 = _RAND_541[20:0];
  _RAND_542 = {1{`RANDOM}};
  way1Tag_29 = _RAND_542[20:0];
  _RAND_543 = {1{`RANDOM}};
  way1Tag_30 = _RAND_543[20:0];
  _RAND_544 = {1{`RANDOM}};
  way1Tag_31 = _RAND_544[20:0];
  _RAND_545 = {1{`RANDOM}};
  way1Tag_32 = _RAND_545[20:0];
  _RAND_546 = {1{`RANDOM}};
  way1Tag_33 = _RAND_546[20:0];
  _RAND_547 = {1{`RANDOM}};
  way1Tag_34 = _RAND_547[20:0];
  _RAND_548 = {1{`RANDOM}};
  way1Tag_35 = _RAND_548[20:0];
  _RAND_549 = {1{`RANDOM}};
  way1Tag_36 = _RAND_549[20:0];
  _RAND_550 = {1{`RANDOM}};
  way1Tag_37 = _RAND_550[20:0];
  _RAND_551 = {1{`RANDOM}};
  way1Tag_38 = _RAND_551[20:0];
  _RAND_552 = {1{`RANDOM}};
  way1Tag_39 = _RAND_552[20:0];
  _RAND_553 = {1{`RANDOM}};
  way1Tag_40 = _RAND_553[20:0];
  _RAND_554 = {1{`RANDOM}};
  way1Tag_41 = _RAND_554[20:0];
  _RAND_555 = {1{`RANDOM}};
  way1Tag_42 = _RAND_555[20:0];
  _RAND_556 = {1{`RANDOM}};
  way1Tag_43 = _RAND_556[20:0];
  _RAND_557 = {1{`RANDOM}};
  way1Tag_44 = _RAND_557[20:0];
  _RAND_558 = {1{`RANDOM}};
  way1Tag_45 = _RAND_558[20:0];
  _RAND_559 = {1{`RANDOM}};
  way1Tag_46 = _RAND_559[20:0];
  _RAND_560 = {1{`RANDOM}};
  way1Tag_47 = _RAND_560[20:0];
  _RAND_561 = {1{`RANDOM}};
  way1Tag_48 = _RAND_561[20:0];
  _RAND_562 = {1{`RANDOM}};
  way1Tag_49 = _RAND_562[20:0];
  _RAND_563 = {1{`RANDOM}};
  way1Tag_50 = _RAND_563[20:0];
  _RAND_564 = {1{`RANDOM}};
  way1Tag_51 = _RAND_564[20:0];
  _RAND_565 = {1{`RANDOM}};
  way1Tag_52 = _RAND_565[20:0];
  _RAND_566 = {1{`RANDOM}};
  way1Tag_53 = _RAND_566[20:0];
  _RAND_567 = {1{`RANDOM}};
  way1Tag_54 = _RAND_567[20:0];
  _RAND_568 = {1{`RANDOM}};
  way1Tag_55 = _RAND_568[20:0];
  _RAND_569 = {1{`RANDOM}};
  way1Tag_56 = _RAND_569[20:0];
  _RAND_570 = {1{`RANDOM}};
  way1Tag_57 = _RAND_570[20:0];
  _RAND_571 = {1{`RANDOM}};
  way1Tag_58 = _RAND_571[20:0];
  _RAND_572 = {1{`RANDOM}};
  way1Tag_59 = _RAND_572[20:0];
  _RAND_573 = {1{`RANDOM}};
  way1Tag_60 = _RAND_573[20:0];
  _RAND_574 = {1{`RANDOM}};
  way1Tag_61 = _RAND_574[20:0];
  _RAND_575 = {1{`RANDOM}};
  way1Tag_62 = _RAND_575[20:0];
  _RAND_576 = {1{`RANDOM}};
  way1Tag_63 = _RAND_576[20:0];
  _RAND_577 = {1{`RANDOM}};
  way1Tag_64 = _RAND_577[20:0];
  _RAND_578 = {1{`RANDOM}};
  way1Tag_65 = _RAND_578[20:0];
  _RAND_579 = {1{`RANDOM}};
  way1Tag_66 = _RAND_579[20:0];
  _RAND_580 = {1{`RANDOM}};
  way1Tag_67 = _RAND_580[20:0];
  _RAND_581 = {1{`RANDOM}};
  way1Tag_68 = _RAND_581[20:0];
  _RAND_582 = {1{`RANDOM}};
  way1Tag_69 = _RAND_582[20:0];
  _RAND_583 = {1{`RANDOM}};
  way1Tag_70 = _RAND_583[20:0];
  _RAND_584 = {1{`RANDOM}};
  way1Tag_71 = _RAND_584[20:0];
  _RAND_585 = {1{`RANDOM}};
  way1Tag_72 = _RAND_585[20:0];
  _RAND_586 = {1{`RANDOM}};
  way1Tag_73 = _RAND_586[20:0];
  _RAND_587 = {1{`RANDOM}};
  way1Tag_74 = _RAND_587[20:0];
  _RAND_588 = {1{`RANDOM}};
  way1Tag_75 = _RAND_588[20:0];
  _RAND_589 = {1{`RANDOM}};
  way1Tag_76 = _RAND_589[20:0];
  _RAND_590 = {1{`RANDOM}};
  way1Tag_77 = _RAND_590[20:0];
  _RAND_591 = {1{`RANDOM}};
  way1Tag_78 = _RAND_591[20:0];
  _RAND_592 = {1{`RANDOM}};
  way1Tag_79 = _RAND_592[20:0];
  _RAND_593 = {1{`RANDOM}};
  way1Tag_80 = _RAND_593[20:0];
  _RAND_594 = {1{`RANDOM}};
  way1Tag_81 = _RAND_594[20:0];
  _RAND_595 = {1{`RANDOM}};
  way1Tag_82 = _RAND_595[20:0];
  _RAND_596 = {1{`RANDOM}};
  way1Tag_83 = _RAND_596[20:0];
  _RAND_597 = {1{`RANDOM}};
  way1Tag_84 = _RAND_597[20:0];
  _RAND_598 = {1{`RANDOM}};
  way1Tag_85 = _RAND_598[20:0];
  _RAND_599 = {1{`RANDOM}};
  way1Tag_86 = _RAND_599[20:0];
  _RAND_600 = {1{`RANDOM}};
  way1Tag_87 = _RAND_600[20:0];
  _RAND_601 = {1{`RANDOM}};
  way1Tag_88 = _RAND_601[20:0];
  _RAND_602 = {1{`RANDOM}};
  way1Tag_89 = _RAND_602[20:0];
  _RAND_603 = {1{`RANDOM}};
  way1Tag_90 = _RAND_603[20:0];
  _RAND_604 = {1{`RANDOM}};
  way1Tag_91 = _RAND_604[20:0];
  _RAND_605 = {1{`RANDOM}};
  way1Tag_92 = _RAND_605[20:0];
  _RAND_606 = {1{`RANDOM}};
  way1Tag_93 = _RAND_606[20:0];
  _RAND_607 = {1{`RANDOM}};
  way1Tag_94 = _RAND_607[20:0];
  _RAND_608 = {1{`RANDOM}};
  way1Tag_95 = _RAND_608[20:0];
  _RAND_609 = {1{`RANDOM}};
  way1Tag_96 = _RAND_609[20:0];
  _RAND_610 = {1{`RANDOM}};
  way1Tag_97 = _RAND_610[20:0];
  _RAND_611 = {1{`RANDOM}};
  way1Tag_98 = _RAND_611[20:0];
  _RAND_612 = {1{`RANDOM}};
  way1Tag_99 = _RAND_612[20:0];
  _RAND_613 = {1{`RANDOM}};
  way1Tag_100 = _RAND_613[20:0];
  _RAND_614 = {1{`RANDOM}};
  way1Tag_101 = _RAND_614[20:0];
  _RAND_615 = {1{`RANDOM}};
  way1Tag_102 = _RAND_615[20:0];
  _RAND_616 = {1{`RANDOM}};
  way1Tag_103 = _RAND_616[20:0];
  _RAND_617 = {1{`RANDOM}};
  way1Tag_104 = _RAND_617[20:0];
  _RAND_618 = {1{`RANDOM}};
  way1Tag_105 = _RAND_618[20:0];
  _RAND_619 = {1{`RANDOM}};
  way1Tag_106 = _RAND_619[20:0];
  _RAND_620 = {1{`RANDOM}};
  way1Tag_107 = _RAND_620[20:0];
  _RAND_621 = {1{`RANDOM}};
  way1Tag_108 = _RAND_621[20:0];
  _RAND_622 = {1{`RANDOM}};
  way1Tag_109 = _RAND_622[20:0];
  _RAND_623 = {1{`RANDOM}};
  way1Tag_110 = _RAND_623[20:0];
  _RAND_624 = {1{`RANDOM}};
  way1Tag_111 = _RAND_624[20:0];
  _RAND_625 = {1{`RANDOM}};
  way1Tag_112 = _RAND_625[20:0];
  _RAND_626 = {1{`RANDOM}};
  way1Tag_113 = _RAND_626[20:0];
  _RAND_627 = {1{`RANDOM}};
  way1Tag_114 = _RAND_627[20:0];
  _RAND_628 = {1{`RANDOM}};
  way1Tag_115 = _RAND_628[20:0];
  _RAND_629 = {1{`RANDOM}};
  way1Tag_116 = _RAND_629[20:0];
  _RAND_630 = {1{`RANDOM}};
  way1Tag_117 = _RAND_630[20:0];
  _RAND_631 = {1{`RANDOM}};
  way1Tag_118 = _RAND_631[20:0];
  _RAND_632 = {1{`RANDOM}};
  way1Tag_119 = _RAND_632[20:0];
  _RAND_633 = {1{`RANDOM}};
  way1Tag_120 = _RAND_633[20:0];
  _RAND_634 = {1{`RANDOM}};
  way1Tag_121 = _RAND_634[20:0];
  _RAND_635 = {1{`RANDOM}};
  way1Tag_122 = _RAND_635[20:0];
  _RAND_636 = {1{`RANDOM}};
  way1Tag_123 = _RAND_636[20:0];
  _RAND_637 = {1{`RANDOM}};
  way1Tag_124 = _RAND_637[20:0];
  _RAND_638 = {1{`RANDOM}};
  way1Tag_125 = _RAND_638[20:0];
  _RAND_639 = {1{`RANDOM}};
  way1Tag_126 = _RAND_639[20:0];
  _RAND_640 = {1{`RANDOM}};
  way1Tag_127 = _RAND_640[20:0];
  _RAND_641 = {1{`RANDOM}};
  way1Age_0 = _RAND_641[0:0];
  _RAND_642 = {1{`RANDOM}};
  way1Age_1 = _RAND_642[0:0];
  _RAND_643 = {1{`RANDOM}};
  way1Age_2 = _RAND_643[0:0];
  _RAND_644 = {1{`RANDOM}};
  way1Age_3 = _RAND_644[0:0];
  _RAND_645 = {1{`RANDOM}};
  way1Age_4 = _RAND_645[0:0];
  _RAND_646 = {1{`RANDOM}};
  way1Age_5 = _RAND_646[0:0];
  _RAND_647 = {1{`RANDOM}};
  way1Age_6 = _RAND_647[0:0];
  _RAND_648 = {1{`RANDOM}};
  way1Age_7 = _RAND_648[0:0];
  _RAND_649 = {1{`RANDOM}};
  way1Age_8 = _RAND_649[0:0];
  _RAND_650 = {1{`RANDOM}};
  way1Age_9 = _RAND_650[0:0];
  _RAND_651 = {1{`RANDOM}};
  way1Age_10 = _RAND_651[0:0];
  _RAND_652 = {1{`RANDOM}};
  way1Age_11 = _RAND_652[0:0];
  _RAND_653 = {1{`RANDOM}};
  way1Age_12 = _RAND_653[0:0];
  _RAND_654 = {1{`RANDOM}};
  way1Age_13 = _RAND_654[0:0];
  _RAND_655 = {1{`RANDOM}};
  way1Age_14 = _RAND_655[0:0];
  _RAND_656 = {1{`RANDOM}};
  way1Age_15 = _RAND_656[0:0];
  _RAND_657 = {1{`RANDOM}};
  way1Age_16 = _RAND_657[0:0];
  _RAND_658 = {1{`RANDOM}};
  way1Age_17 = _RAND_658[0:0];
  _RAND_659 = {1{`RANDOM}};
  way1Age_18 = _RAND_659[0:0];
  _RAND_660 = {1{`RANDOM}};
  way1Age_19 = _RAND_660[0:0];
  _RAND_661 = {1{`RANDOM}};
  way1Age_20 = _RAND_661[0:0];
  _RAND_662 = {1{`RANDOM}};
  way1Age_21 = _RAND_662[0:0];
  _RAND_663 = {1{`RANDOM}};
  way1Age_22 = _RAND_663[0:0];
  _RAND_664 = {1{`RANDOM}};
  way1Age_23 = _RAND_664[0:0];
  _RAND_665 = {1{`RANDOM}};
  way1Age_24 = _RAND_665[0:0];
  _RAND_666 = {1{`RANDOM}};
  way1Age_25 = _RAND_666[0:0];
  _RAND_667 = {1{`RANDOM}};
  way1Age_26 = _RAND_667[0:0];
  _RAND_668 = {1{`RANDOM}};
  way1Age_27 = _RAND_668[0:0];
  _RAND_669 = {1{`RANDOM}};
  way1Age_28 = _RAND_669[0:0];
  _RAND_670 = {1{`RANDOM}};
  way1Age_29 = _RAND_670[0:0];
  _RAND_671 = {1{`RANDOM}};
  way1Age_30 = _RAND_671[0:0];
  _RAND_672 = {1{`RANDOM}};
  way1Age_31 = _RAND_672[0:0];
  _RAND_673 = {1{`RANDOM}};
  way1Age_32 = _RAND_673[0:0];
  _RAND_674 = {1{`RANDOM}};
  way1Age_33 = _RAND_674[0:0];
  _RAND_675 = {1{`RANDOM}};
  way1Age_34 = _RAND_675[0:0];
  _RAND_676 = {1{`RANDOM}};
  way1Age_35 = _RAND_676[0:0];
  _RAND_677 = {1{`RANDOM}};
  way1Age_36 = _RAND_677[0:0];
  _RAND_678 = {1{`RANDOM}};
  way1Age_37 = _RAND_678[0:0];
  _RAND_679 = {1{`RANDOM}};
  way1Age_38 = _RAND_679[0:0];
  _RAND_680 = {1{`RANDOM}};
  way1Age_39 = _RAND_680[0:0];
  _RAND_681 = {1{`RANDOM}};
  way1Age_40 = _RAND_681[0:0];
  _RAND_682 = {1{`RANDOM}};
  way1Age_41 = _RAND_682[0:0];
  _RAND_683 = {1{`RANDOM}};
  way1Age_42 = _RAND_683[0:0];
  _RAND_684 = {1{`RANDOM}};
  way1Age_43 = _RAND_684[0:0];
  _RAND_685 = {1{`RANDOM}};
  way1Age_44 = _RAND_685[0:0];
  _RAND_686 = {1{`RANDOM}};
  way1Age_45 = _RAND_686[0:0];
  _RAND_687 = {1{`RANDOM}};
  way1Age_46 = _RAND_687[0:0];
  _RAND_688 = {1{`RANDOM}};
  way1Age_47 = _RAND_688[0:0];
  _RAND_689 = {1{`RANDOM}};
  way1Age_48 = _RAND_689[0:0];
  _RAND_690 = {1{`RANDOM}};
  way1Age_49 = _RAND_690[0:0];
  _RAND_691 = {1{`RANDOM}};
  way1Age_50 = _RAND_691[0:0];
  _RAND_692 = {1{`RANDOM}};
  way1Age_51 = _RAND_692[0:0];
  _RAND_693 = {1{`RANDOM}};
  way1Age_52 = _RAND_693[0:0];
  _RAND_694 = {1{`RANDOM}};
  way1Age_53 = _RAND_694[0:0];
  _RAND_695 = {1{`RANDOM}};
  way1Age_54 = _RAND_695[0:0];
  _RAND_696 = {1{`RANDOM}};
  way1Age_55 = _RAND_696[0:0];
  _RAND_697 = {1{`RANDOM}};
  way1Age_56 = _RAND_697[0:0];
  _RAND_698 = {1{`RANDOM}};
  way1Age_57 = _RAND_698[0:0];
  _RAND_699 = {1{`RANDOM}};
  way1Age_58 = _RAND_699[0:0];
  _RAND_700 = {1{`RANDOM}};
  way1Age_59 = _RAND_700[0:0];
  _RAND_701 = {1{`RANDOM}};
  way1Age_60 = _RAND_701[0:0];
  _RAND_702 = {1{`RANDOM}};
  way1Age_61 = _RAND_702[0:0];
  _RAND_703 = {1{`RANDOM}};
  way1Age_62 = _RAND_703[0:0];
  _RAND_704 = {1{`RANDOM}};
  way1Age_63 = _RAND_704[0:0];
  _RAND_705 = {1{`RANDOM}};
  way1Age_64 = _RAND_705[0:0];
  _RAND_706 = {1{`RANDOM}};
  way1Age_65 = _RAND_706[0:0];
  _RAND_707 = {1{`RANDOM}};
  way1Age_66 = _RAND_707[0:0];
  _RAND_708 = {1{`RANDOM}};
  way1Age_67 = _RAND_708[0:0];
  _RAND_709 = {1{`RANDOM}};
  way1Age_68 = _RAND_709[0:0];
  _RAND_710 = {1{`RANDOM}};
  way1Age_69 = _RAND_710[0:0];
  _RAND_711 = {1{`RANDOM}};
  way1Age_70 = _RAND_711[0:0];
  _RAND_712 = {1{`RANDOM}};
  way1Age_71 = _RAND_712[0:0];
  _RAND_713 = {1{`RANDOM}};
  way1Age_72 = _RAND_713[0:0];
  _RAND_714 = {1{`RANDOM}};
  way1Age_73 = _RAND_714[0:0];
  _RAND_715 = {1{`RANDOM}};
  way1Age_74 = _RAND_715[0:0];
  _RAND_716 = {1{`RANDOM}};
  way1Age_75 = _RAND_716[0:0];
  _RAND_717 = {1{`RANDOM}};
  way1Age_76 = _RAND_717[0:0];
  _RAND_718 = {1{`RANDOM}};
  way1Age_77 = _RAND_718[0:0];
  _RAND_719 = {1{`RANDOM}};
  way1Age_78 = _RAND_719[0:0];
  _RAND_720 = {1{`RANDOM}};
  way1Age_79 = _RAND_720[0:0];
  _RAND_721 = {1{`RANDOM}};
  way1Age_80 = _RAND_721[0:0];
  _RAND_722 = {1{`RANDOM}};
  way1Age_81 = _RAND_722[0:0];
  _RAND_723 = {1{`RANDOM}};
  way1Age_82 = _RAND_723[0:0];
  _RAND_724 = {1{`RANDOM}};
  way1Age_83 = _RAND_724[0:0];
  _RAND_725 = {1{`RANDOM}};
  way1Age_84 = _RAND_725[0:0];
  _RAND_726 = {1{`RANDOM}};
  way1Age_85 = _RAND_726[0:0];
  _RAND_727 = {1{`RANDOM}};
  way1Age_86 = _RAND_727[0:0];
  _RAND_728 = {1{`RANDOM}};
  way1Age_87 = _RAND_728[0:0];
  _RAND_729 = {1{`RANDOM}};
  way1Age_88 = _RAND_729[0:0];
  _RAND_730 = {1{`RANDOM}};
  way1Age_89 = _RAND_730[0:0];
  _RAND_731 = {1{`RANDOM}};
  way1Age_90 = _RAND_731[0:0];
  _RAND_732 = {1{`RANDOM}};
  way1Age_91 = _RAND_732[0:0];
  _RAND_733 = {1{`RANDOM}};
  way1Age_92 = _RAND_733[0:0];
  _RAND_734 = {1{`RANDOM}};
  way1Age_93 = _RAND_734[0:0];
  _RAND_735 = {1{`RANDOM}};
  way1Age_94 = _RAND_735[0:0];
  _RAND_736 = {1{`RANDOM}};
  way1Age_95 = _RAND_736[0:0];
  _RAND_737 = {1{`RANDOM}};
  way1Age_96 = _RAND_737[0:0];
  _RAND_738 = {1{`RANDOM}};
  way1Age_97 = _RAND_738[0:0];
  _RAND_739 = {1{`RANDOM}};
  way1Age_98 = _RAND_739[0:0];
  _RAND_740 = {1{`RANDOM}};
  way1Age_99 = _RAND_740[0:0];
  _RAND_741 = {1{`RANDOM}};
  way1Age_100 = _RAND_741[0:0];
  _RAND_742 = {1{`RANDOM}};
  way1Age_101 = _RAND_742[0:0];
  _RAND_743 = {1{`RANDOM}};
  way1Age_102 = _RAND_743[0:0];
  _RAND_744 = {1{`RANDOM}};
  way1Age_103 = _RAND_744[0:0];
  _RAND_745 = {1{`RANDOM}};
  way1Age_104 = _RAND_745[0:0];
  _RAND_746 = {1{`RANDOM}};
  way1Age_105 = _RAND_746[0:0];
  _RAND_747 = {1{`RANDOM}};
  way1Age_106 = _RAND_747[0:0];
  _RAND_748 = {1{`RANDOM}};
  way1Age_107 = _RAND_748[0:0];
  _RAND_749 = {1{`RANDOM}};
  way1Age_108 = _RAND_749[0:0];
  _RAND_750 = {1{`RANDOM}};
  way1Age_109 = _RAND_750[0:0];
  _RAND_751 = {1{`RANDOM}};
  way1Age_110 = _RAND_751[0:0];
  _RAND_752 = {1{`RANDOM}};
  way1Age_111 = _RAND_752[0:0];
  _RAND_753 = {1{`RANDOM}};
  way1Age_112 = _RAND_753[0:0];
  _RAND_754 = {1{`RANDOM}};
  way1Age_113 = _RAND_754[0:0];
  _RAND_755 = {1{`RANDOM}};
  way1Age_114 = _RAND_755[0:0];
  _RAND_756 = {1{`RANDOM}};
  way1Age_115 = _RAND_756[0:0];
  _RAND_757 = {1{`RANDOM}};
  way1Age_116 = _RAND_757[0:0];
  _RAND_758 = {1{`RANDOM}};
  way1Age_117 = _RAND_758[0:0];
  _RAND_759 = {1{`RANDOM}};
  way1Age_118 = _RAND_759[0:0];
  _RAND_760 = {1{`RANDOM}};
  way1Age_119 = _RAND_760[0:0];
  _RAND_761 = {1{`RANDOM}};
  way1Age_120 = _RAND_761[0:0];
  _RAND_762 = {1{`RANDOM}};
  way1Age_121 = _RAND_762[0:0];
  _RAND_763 = {1{`RANDOM}};
  way1Age_122 = _RAND_763[0:0];
  _RAND_764 = {1{`RANDOM}};
  way1Age_123 = _RAND_764[0:0];
  _RAND_765 = {1{`RANDOM}};
  way1Age_124 = _RAND_765[0:0];
  _RAND_766 = {1{`RANDOM}};
  way1Age_125 = _RAND_766[0:0];
  _RAND_767 = {1{`RANDOM}};
  way1Age_126 = _RAND_767[0:0];
  _RAND_768 = {1{`RANDOM}};
  way1Age_127 = _RAND_768[0:0];
  _RAND_769 = {1{`RANDOM}};
  state = _RAND_769[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module DCache(
  input          clock,
  input          reset,
  input          io_dmem_data_valid,
  output         io_dmem_data_ready,
  input          io_dmem_data_req,
  input  [31:0]  io_dmem_data_addr,
  input  [1:0]   io_dmem_data_size,
  input  [7:0]   io_dmem_data_strb,
  output [63:0]  io_dmem_data_read,
  input  [127:0] io_dmem_data_write,
  output         io_out_data_valid,
  input          io_out_data_ready,
  output         io_out_data_req,
  output [31:0]  io_out_data_addr,
  output [7:0]   io_out_data_strb,
  input  [127:0] io_out_data_read,
  output [127:0] io_out_data_write
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_645;
  reg [31:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_649;
  reg [31:0] _RAND_650;
  reg [31:0] _RAND_651;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
  reg [31:0] _RAND_654;
  reg [31:0] _RAND_655;
  reg [31:0] _RAND_656;
  reg [31:0] _RAND_657;
  reg [31:0] _RAND_658;
  reg [31:0] _RAND_659;
  reg [31:0] _RAND_660;
  reg [31:0] _RAND_661;
  reg [31:0] _RAND_662;
  reg [31:0] _RAND_663;
  reg [31:0] _RAND_664;
  reg [31:0] _RAND_665;
  reg [31:0] _RAND_666;
  reg [31:0] _RAND_667;
  reg [31:0] _RAND_668;
  reg [31:0] _RAND_669;
  reg [31:0] _RAND_670;
  reg [31:0] _RAND_671;
  reg [31:0] _RAND_672;
  reg [31:0] _RAND_673;
  reg [31:0] _RAND_674;
  reg [31:0] _RAND_675;
  reg [31:0] _RAND_676;
  reg [31:0] _RAND_677;
  reg [31:0] _RAND_678;
  reg [31:0] _RAND_679;
  reg [31:0] _RAND_680;
  reg [31:0] _RAND_681;
  reg [31:0] _RAND_682;
  reg [31:0] _RAND_683;
  reg [31:0] _RAND_684;
  reg [31:0] _RAND_685;
  reg [31:0] _RAND_686;
  reg [31:0] _RAND_687;
  reg [31:0] _RAND_688;
  reg [31:0] _RAND_689;
  reg [31:0] _RAND_690;
  reg [31:0] _RAND_691;
  reg [31:0] _RAND_692;
  reg [31:0] _RAND_693;
  reg [31:0] _RAND_694;
  reg [31:0] _RAND_695;
  reg [31:0] _RAND_696;
  reg [31:0] _RAND_697;
  reg [31:0] _RAND_698;
  reg [31:0] _RAND_699;
  reg [31:0] _RAND_700;
  reg [31:0] _RAND_701;
  reg [31:0] _RAND_702;
  reg [31:0] _RAND_703;
  reg [31:0] _RAND_704;
  reg [31:0] _RAND_705;
  reg [31:0] _RAND_706;
  reg [31:0] _RAND_707;
  reg [31:0] _RAND_708;
  reg [31:0] _RAND_709;
  reg [31:0] _RAND_710;
  reg [31:0] _RAND_711;
  reg [31:0] _RAND_712;
  reg [31:0] _RAND_713;
  reg [31:0] _RAND_714;
  reg [31:0] _RAND_715;
  reg [31:0] _RAND_716;
  reg [31:0] _RAND_717;
  reg [31:0] _RAND_718;
  reg [31:0] _RAND_719;
  reg [31:0] _RAND_720;
  reg [31:0] _RAND_721;
  reg [31:0] _RAND_722;
  reg [31:0] _RAND_723;
  reg [31:0] _RAND_724;
  reg [31:0] _RAND_725;
  reg [31:0] _RAND_726;
  reg [31:0] _RAND_727;
  reg [31:0] _RAND_728;
  reg [31:0] _RAND_729;
  reg [31:0] _RAND_730;
  reg [31:0] _RAND_731;
  reg [31:0] _RAND_732;
  reg [31:0] _RAND_733;
  reg [31:0] _RAND_734;
  reg [31:0] _RAND_735;
  reg [31:0] _RAND_736;
  reg [31:0] _RAND_737;
  reg [31:0] _RAND_738;
  reg [31:0] _RAND_739;
  reg [31:0] _RAND_740;
  reg [31:0] _RAND_741;
  reg [31:0] _RAND_742;
  reg [31:0] _RAND_743;
  reg [31:0] _RAND_744;
  reg [31:0] _RAND_745;
  reg [31:0] _RAND_746;
  reg [31:0] _RAND_747;
  reg [31:0] _RAND_748;
  reg [31:0] _RAND_749;
  reg [31:0] _RAND_750;
  reg [31:0] _RAND_751;
  reg [31:0] _RAND_752;
  reg [31:0] _RAND_753;
  reg [31:0] _RAND_754;
  reg [31:0] _RAND_755;
  reg [31:0] _RAND_756;
  reg [31:0] _RAND_757;
  reg [31:0] _RAND_758;
  reg [31:0] _RAND_759;
  reg [31:0] _RAND_760;
  reg [31:0] _RAND_761;
  reg [31:0] _RAND_762;
  reg [31:0] _RAND_763;
  reg [31:0] _RAND_764;
  reg [31:0] _RAND_765;
  reg [31:0] _RAND_766;
  reg [31:0] _RAND_767;
  reg [31:0] _RAND_768;
  reg [31:0] _RAND_769;
  reg [31:0] _RAND_770;
  reg [31:0] _RAND_771;
  reg [31:0] _RAND_772;
  reg [31:0] _RAND_773;
  reg [31:0] _RAND_774;
  reg [31:0] _RAND_775;
  reg [31:0] _RAND_776;
  reg [31:0] _RAND_777;
  reg [31:0] _RAND_778;
  reg [31:0] _RAND_779;
  reg [31:0] _RAND_780;
  reg [31:0] _RAND_781;
  reg [31:0] _RAND_782;
  reg [31:0] _RAND_783;
  reg [31:0] _RAND_784;
  reg [31:0] _RAND_785;
  reg [31:0] _RAND_786;
  reg [31:0] _RAND_787;
  reg [31:0] _RAND_788;
  reg [31:0] _RAND_789;
  reg [31:0] _RAND_790;
  reg [31:0] _RAND_791;
  reg [31:0] _RAND_792;
  reg [31:0] _RAND_793;
  reg [31:0] _RAND_794;
  reg [31:0] _RAND_795;
  reg [31:0] _RAND_796;
  reg [31:0] _RAND_797;
  reg [31:0] _RAND_798;
  reg [31:0] _RAND_799;
  reg [31:0] _RAND_800;
  reg [31:0] _RAND_801;
  reg [31:0] _RAND_802;
  reg [31:0] _RAND_803;
  reg [31:0] _RAND_804;
  reg [31:0] _RAND_805;
  reg [31:0] _RAND_806;
  reg [31:0] _RAND_807;
  reg [31:0] _RAND_808;
  reg [31:0] _RAND_809;
  reg [31:0] _RAND_810;
  reg [31:0] _RAND_811;
  reg [31:0] _RAND_812;
  reg [31:0] _RAND_813;
  reg [31:0] _RAND_814;
  reg [31:0] _RAND_815;
  reg [31:0] _RAND_816;
  reg [31:0] _RAND_817;
  reg [31:0] _RAND_818;
  reg [31:0] _RAND_819;
  reg [31:0] _RAND_820;
  reg [31:0] _RAND_821;
  reg [31:0] _RAND_822;
  reg [31:0] _RAND_823;
  reg [31:0] _RAND_824;
  reg [31:0] _RAND_825;
  reg [31:0] _RAND_826;
  reg [31:0] _RAND_827;
  reg [31:0] _RAND_828;
  reg [31:0] _RAND_829;
  reg [31:0] _RAND_830;
  reg [31:0] _RAND_831;
  reg [31:0] _RAND_832;
  reg [31:0] _RAND_833;
  reg [31:0] _RAND_834;
  reg [31:0] _RAND_835;
  reg [31:0] _RAND_836;
  reg [31:0] _RAND_837;
  reg [31:0] _RAND_838;
  reg [31:0] _RAND_839;
  reg [31:0] _RAND_840;
  reg [31:0] _RAND_841;
  reg [31:0] _RAND_842;
  reg [31:0] _RAND_843;
  reg [31:0] _RAND_844;
  reg [31:0] _RAND_845;
  reg [31:0] _RAND_846;
  reg [31:0] _RAND_847;
  reg [31:0] _RAND_848;
  reg [31:0] _RAND_849;
  reg [31:0] _RAND_850;
  reg [31:0] _RAND_851;
  reg [31:0] _RAND_852;
  reg [31:0] _RAND_853;
  reg [31:0] _RAND_854;
  reg [31:0] _RAND_855;
  reg [31:0] _RAND_856;
  reg [31:0] _RAND_857;
  reg [31:0] _RAND_858;
  reg [31:0] _RAND_859;
  reg [31:0] _RAND_860;
  reg [31:0] _RAND_861;
  reg [31:0] _RAND_862;
  reg [31:0] _RAND_863;
  reg [31:0] _RAND_864;
  reg [31:0] _RAND_865;
  reg [31:0] _RAND_866;
  reg [31:0] _RAND_867;
  reg [31:0] _RAND_868;
  reg [31:0] _RAND_869;
  reg [31:0] _RAND_870;
  reg [31:0] _RAND_871;
  reg [31:0] _RAND_872;
  reg [31:0] _RAND_873;
  reg [31:0] _RAND_874;
  reg [31:0] _RAND_875;
  reg [31:0] _RAND_876;
  reg [31:0] _RAND_877;
  reg [31:0] _RAND_878;
  reg [31:0] _RAND_879;
  reg [31:0] _RAND_880;
  reg [31:0] _RAND_881;
  reg [31:0] _RAND_882;
  reg [31:0] _RAND_883;
  reg [31:0] _RAND_884;
  reg [31:0] _RAND_885;
  reg [31:0] _RAND_886;
  reg [31:0] _RAND_887;
  reg [31:0] _RAND_888;
  reg [31:0] _RAND_889;
  reg [31:0] _RAND_890;
  reg [31:0] _RAND_891;
  reg [31:0] _RAND_892;
  reg [31:0] _RAND_893;
  reg [31:0] _RAND_894;
  reg [31:0] _RAND_895;
  reg [31:0] _RAND_896;
  reg [31:0] _RAND_897;
  reg [31:0] _RAND_898;
  reg [31:0] _RAND_899;
  reg [31:0] _RAND_900;
  reg [31:0] _RAND_901;
  reg [31:0] _RAND_902;
  reg [31:0] _RAND_903;
  reg [31:0] _RAND_904;
  reg [31:0] _RAND_905;
  reg [31:0] _RAND_906;
  reg [31:0] _RAND_907;
  reg [31:0] _RAND_908;
  reg [31:0] _RAND_909;
  reg [31:0] _RAND_910;
  reg [31:0] _RAND_911;
  reg [31:0] _RAND_912;
  reg [31:0] _RAND_913;
  reg [31:0] _RAND_914;
  reg [31:0] _RAND_915;
  reg [31:0] _RAND_916;
  reg [31:0] _RAND_917;
  reg [31:0] _RAND_918;
  reg [31:0] _RAND_919;
  reg [31:0] _RAND_920;
  reg [31:0] _RAND_921;
  reg [31:0] _RAND_922;
  reg [31:0] _RAND_923;
  reg [31:0] _RAND_924;
  reg [31:0] _RAND_925;
  reg [31:0] _RAND_926;
  reg [31:0] _RAND_927;
  reg [31:0] _RAND_928;
  reg [31:0] _RAND_929;
  reg [31:0] _RAND_930;
  reg [31:0] _RAND_931;
  reg [31:0] _RAND_932;
  reg [31:0] _RAND_933;
  reg [31:0] _RAND_934;
  reg [31:0] _RAND_935;
  reg [31:0] _RAND_936;
  reg [31:0] _RAND_937;
  reg [31:0] _RAND_938;
  reg [31:0] _RAND_939;
  reg [31:0] _RAND_940;
  reg [31:0] _RAND_941;
  reg [31:0] _RAND_942;
  reg [31:0] _RAND_943;
  reg [31:0] _RAND_944;
  reg [31:0] _RAND_945;
  reg [31:0] _RAND_946;
  reg [31:0] _RAND_947;
  reg [31:0] _RAND_948;
  reg [31:0] _RAND_949;
  reg [31:0] _RAND_950;
  reg [31:0] _RAND_951;
  reg [31:0] _RAND_952;
  reg [31:0] _RAND_953;
  reg [31:0] _RAND_954;
  reg [31:0] _RAND_955;
  reg [31:0] _RAND_956;
  reg [31:0] _RAND_957;
  reg [31:0] _RAND_958;
  reg [31:0] _RAND_959;
  reg [31:0] _RAND_960;
  reg [31:0] _RAND_961;
  reg [31:0] _RAND_962;
  reg [31:0] _RAND_963;
  reg [31:0] _RAND_964;
  reg [31:0] _RAND_965;
  reg [31:0] _RAND_966;
  reg [31:0] _RAND_967;
  reg [31:0] _RAND_968;
  reg [31:0] _RAND_969;
  reg [31:0] _RAND_970;
  reg [31:0] _RAND_971;
  reg [31:0] _RAND_972;
  reg [31:0] _RAND_973;
  reg [31:0] _RAND_974;
  reg [31:0] _RAND_975;
  reg [31:0] _RAND_976;
  reg [31:0] _RAND_977;
  reg [31:0] _RAND_978;
  reg [31:0] _RAND_979;
  reg [31:0] _RAND_980;
  reg [31:0] _RAND_981;
  reg [31:0] _RAND_982;
  reg [31:0] _RAND_983;
  reg [31:0] _RAND_984;
  reg [31:0] _RAND_985;
  reg [31:0] _RAND_986;
  reg [31:0] _RAND_987;
  reg [31:0] _RAND_988;
  reg [31:0] _RAND_989;
  reg [31:0] _RAND_990;
  reg [31:0] _RAND_991;
  reg [31:0] _RAND_992;
  reg [31:0] _RAND_993;
  reg [31:0] _RAND_994;
  reg [31:0] _RAND_995;
  reg [31:0] _RAND_996;
  reg [31:0] _RAND_997;
  reg [31:0] _RAND_998;
  reg [31:0] _RAND_999;
  reg [31:0] _RAND_1000;
  reg [31:0] _RAND_1001;
  reg [31:0] _RAND_1002;
  reg [31:0] _RAND_1003;
  reg [31:0] _RAND_1004;
  reg [31:0] _RAND_1005;
  reg [31:0] _RAND_1006;
  reg [31:0] _RAND_1007;
  reg [31:0] _RAND_1008;
  reg [31:0] _RAND_1009;
  reg [31:0] _RAND_1010;
  reg [31:0] _RAND_1011;
  reg [31:0] _RAND_1012;
  reg [31:0] _RAND_1013;
  reg [31:0] _RAND_1014;
  reg [31:0] _RAND_1015;
  reg [31:0] _RAND_1016;
  reg [31:0] _RAND_1017;
  reg [31:0] _RAND_1018;
  reg [31:0] _RAND_1019;
  reg [31:0] _RAND_1020;
  reg [31:0] _RAND_1021;
  reg [31:0] _RAND_1022;
  reg [31:0] _RAND_1023;
  reg [31:0] _RAND_1024;
  reg [31:0] _RAND_1025;
`endif // RANDOMIZE_REG_INIT
  wire [127:0] req_Q; // @[DCache.scala 253:19]
  wire  req_CLK; // @[DCache.scala 253:19]
  wire  req_CEN; // @[DCache.scala 253:19]
  wire  req_WEN; // @[DCache.scala 253:19]
  wire [127:0] req_BWEN; // @[DCache.scala 253:19]
  wire [7:0] req_A; // @[DCache.scala 253:19]
  wire [127:0] req_D; // @[DCache.scala 253:19]
  reg  way0V_0; // @[DCache.scala 33:26]
  reg  way0V_1; // @[DCache.scala 33:26]
  reg  way0V_2; // @[DCache.scala 33:26]
  reg  way0V_3; // @[DCache.scala 33:26]
  reg  way0V_4; // @[DCache.scala 33:26]
  reg  way0V_5; // @[DCache.scala 33:26]
  reg  way0V_6; // @[DCache.scala 33:26]
  reg  way0V_7; // @[DCache.scala 33:26]
  reg  way0V_8; // @[DCache.scala 33:26]
  reg  way0V_9; // @[DCache.scala 33:26]
  reg  way0V_10; // @[DCache.scala 33:26]
  reg  way0V_11; // @[DCache.scala 33:26]
  reg  way0V_12; // @[DCache.scala 33:26]
  reg  way0V_13; // @[DCache.scala 33:26]
  reg  way0V_14; // @[DCache.scala 33:26]
  reg  way0V_15; // @[DCache.scala 33:26]
  reg  way0V_16; // @[DCache.scala 33:26]
  reg  way0V_17; // @[DCache.scala 33:26]
  reg  way0V_18; // @[DCache.scala 33:26]
  reg  way0V_19; // @[DCache.scala 33:26]
  reg  way0V_20; // @[DCache.scala 33:26]
  reg  way0V_21; // @[DCache.scala 33:26]
  reg  way0V_22; // @[DCache.scala 33:26]
  reg  way0V_23; // @[DCache.scala 33:26]
  reg  way0V_24; // @[DCache.scala 33:26]
  reg  way0V_25; // @[DCache.scala 33:26]
  reg  way0V_26; // @[DCache.scala 33:26]
  reg  way0V_27; // @[DCache.scala 33:26]
  reg  way0V_28; // @[DCache.scala 33:26]
  reg  way0V_29; // @[DCache.scala 33:26]
  reg  way0V_30; // @[DCache.scala 33:26]
  reg  way0V_31; // @[DCache.scala 33:26]
  reg  way0V_32; // @[DCache.scala 33:26]
  reg  way0V_33; // @[DCache.scala 33:26]
  reg  way0V_34; // @[DCache.scala 33:26]
  reg  way0V_35; // @[DCache.scala 33:26]
  reg  way0V_36; // @[DCache.scala 33:26]
  reg  way0V_37; // @[DCache.scala 33:26]
  reg  way0V_38; // @[DCache.scala 33:26]
  reg  way0V_39; // @[DCache.scala 33:26]
  reg  way0V_40; // @[DCache.scala 33:26]
  reg  way0V_41; // @[DCache.scala 33:26]
  reg  way0V_42; // @[DCache.scala 33:26]
  reg  way0V_43; // @[DCache.scala 33:26]
  reg  way0V_44; // @[DCache.scala 33:26]
  reg  way0V_45; // @[DCache.scala 33:26]
  reg  way0V_46; // @[DCache.scala 33:26]
  reg  way0V_47; // @[DCache.scala 33:26]
  reg  way0V_48; // @[DCache.scala 33:26]
  reg  way0V_49; // @[DCache.scala 33:26]
  reg  way0V_50; // @[DCache.scala 33:26]
  reg  way0V_51; // @[DCache.scala 33:26]
  reg  way0V_52; // @[DCache.scala 33:26]
  reg  way0V_53; // @[DCache.scala 33:26]
  reg  way0V_54; // @[DCache.scala 33:26]
  reg  way0V_55; // @[DCache.scala 33:26]
  reg  way0V_56; // @[DCache.scala 33:26]
  reg  way0V_57; // @[DCache.scala 33:26]
  reg  way0V_58; // @[DCache.scala 33:26]
  reg  way0V_59; // @[DCache.scala 33:26]
  reg  way0V_60; // @[DCache.scala 33:26]
  reg  way0V_61; // @[DCache.scala 33:26]
  reg  way0V_62; // @[DCache.scala 33:26]
  reg  way0V_63; // @[DCache.scala 33:26]
  reg  way0V_64; // @[DCache.scala 33:26]
  reg  way0V_65; // @[DCache.scala 33:26]
  reg  way0V_66; // @[DCache.scala 33:26]
  reg  way0V_67; // @[DCache.scala 33:26]
  reg  way0V_68; // @[DCache.scala 33:26]
  reg  way0V_69; // @[DCache.scala 33:26]
  reg  way0V_70; // @[DCache.scala 33:26]
  reg  way0V_71; // @[DCache.scala 33:26]
  reg  way0V_72; // @[DCache.scala 33:26]
  reg  way0V_73; // @[DCache.scala 33:26]
  reg  way0V_74; // @[DCache.scala 33:26]
  reg  way0V_75; // @[DCache.scala 33:26]
  reg  way0V_76; // @[DCache.scala 33:26]
  reg  way0V_77; // @[DCache.scala 33:26]
  reg  way0V_78; // @[DCache.scala 33:26]
  reg  way0V_79; // @[DCache.scala 33:26]
  reg  way0V_80; // @[DCache.scala 33:26]
  reg  way0V_81; // @[DCache.scala 33:26]
  reg  way0V_82; // @[DCache.scala 33:26]
  reg  way0V_83; // @[DCache.scala 33:26]
  reg  way0V_84; // @[DCache.scala 33:26]
  reg  way0V_85; // @[DCache.scala 33:26]
  reg  way0V_86; // @[DCache.scala 33:26]
  reg  way0V_87; // @[DCache.scala 33:26]
  reg  way0V_88; // @[DCache.scala 33:26]
  reg  way0V_89; // @[DCache.scala 33:26]
  reg  way0V_90; // @[DCache.scala 33:26]
  reg  way0V_91; // @[DCache.scala 33:26]
  reg  way0V_92; // @[DCache.scala 33:26]
  reg  way0V_93; // @[DCache.scala 33:26]
  reg  way0V_94; // @[DCache.scala 33:26]
  reg  way0V_95; // @[DCache.scala 33:26]
  reg  way0V_96; // @[DCache.scala 33:26]
  reg  way0V_97; // @[DCache.scala 33:26]
  reg  way0V_98; // @[DCache.scala 33:26]
  reg  way0V_99; // @[DCache.scala 33:26]
  reg  way0V_100; // @[DCache.scala 33:26]
  reg  way0V_101; // @[DCache.scala 33:26]
  reg  way0V_102; // @[DCache.scala 33:26]
  reg  way0V_103; // @[DCache.scala 33:26]
  reg  way0V_104; // @[DCache.scala 33:26]
  reg  way0V_105; // @[DCache.scala 33:26]
  reg  way0V_106; // @[DCache.scala 33:26]
  reg  way0V_107; // @[DCache.scala 33:26]
  reg  way0V_108; // @[DCache.scala 33:26]
  reg  way0V_109; // @[DCache.scala 33:26]
  reg  way0V_110; // @[DCache.scala 33:26]
  reg  way0V_111; // @[DCache.scala 33:26]
  reg  way0V_112; // @[DCache.scala 33:26]
  reg  way0V_113; // @[DCache.scala 33:26]
  reg  way0V_114; // @[DCache.scala 33:26]
  reg  way0V_115; // @[DCache.scala 33:26]
  reg  way0V_116; // @[DCache.scala 33:26]
  reg  way0V_117; // @[DCache.scala 33:26]
  reg  way0V_118; // @[DCache.scala 33:26]
  reg  way0V_119; // @[DCache.scala 33:26]
  reg  way0V_120; // @[DCache.scala 33:26]
  reg  way0V_121; // @[DCache.scala 33:26]
  reg  way0V_122; // @[DCache.scala 33:26]
  reg  way0V_123; // @[DCache.scala 33:26]
  reg  way0V_124; // @[DCache.scala 33:26]
  reg  way0V_125; // @[DCache.scala 33:26]
  reg  way0V_126; // @[DCache.scala 33:26]
  reg  way0V_127; // @[DCache.scala 33:26]
  reg [20:0] way0Tag_0; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_1; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_2; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_3; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_4; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_5; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_6; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_7; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_8; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_9; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_10; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_11; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_12; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_13; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_14; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_15; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_16; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_17; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_18; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_19; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_20; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_21; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_22; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_23; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_24; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_25; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_26; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_27; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_28; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_29; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_30; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_31; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_32; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_33; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_34; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_35; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_36; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_37; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_38; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_39; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_40; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_41; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_42; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_43; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_44; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_45; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_46; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_47; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_48; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_49; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_50; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_51; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_52; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_53; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_54; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_55; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_56; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_57; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_58; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_59; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_60; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_61; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_62; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_63; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_64; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_65; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_66; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_67; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_68; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_69; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_70; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_71; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_72; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_73; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_74; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_75; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_76; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_77; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_78; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_79; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_80; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_81; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_82; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_83; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_84; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_85; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_86; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_87; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_88; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_89; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_90; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_91; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_92; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_93; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_94; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_95; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_96; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_97; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_98; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_99; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_100; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_101; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_102; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_103; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_104; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_105; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_106; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_107; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_108; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_109; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_110; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_111; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_112; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_113; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_114; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_115; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_116; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_117; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_118; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_119; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_120; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_121; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_122; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_123; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_124; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_125; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_126; // @[DCache.scala 34:26]
  reg [20:0] way0Tag_127; // @[DCache.scala 34:26]
  reg  way0Age_0; // @[DCache.scala 36:26]
  reg  way0Age_1; // @[DCache.scala 36:26]
  reg  way0Age_2; // @[DCache.scala 36:26]
  reg  way0Age_3; // @[DCache.scala 36:26]
  reg  way0Age_4; // @[DCache.scala 36:26]
  reg  way0Age_5; // @[DCache.scala 36:26]
  reg  way0Age_6; // @[DCache.scala 36:26]
  reg  way0Age_7; // @[DCache.scala 36:26]
  reg  way0Age_8; // @[DCache.scala 36:26]
  reg  way0Age_9; // @[DCache.scala 36:26]
  reg  way0Age_10; // @[DCache.scala 36:26]
  reg  way0Age_11; // @[DCache.scala 36:26]
  reg  way0Age_12; // @[DCache.scala 36:26]
  reg  way0Age_13; // @[DCache.scala 36:26]
  reg  way0Age_14; // @[DCache.scala 36:26]
  reg  way0Age_15; // @[DCache.scala 36:26]
  reg  way0Age_16; // @[DCache.scala 36:26]
  reg  way0Age_17; // @[DCache.scala 36:26]
  reg  way0Age_18; // @[DCache.scala 36:26]
  reg  way0Age_19; // @[DCache.scala 36:26]
  reg  way0Age_20; // @[DCache.scala 36:26]
  reg  way0Age_21; // @[DCache.scala 36:26]
  reg  way0Age_22; // @[DCache.scala 36:26]
  reg  way0Age_23; // @[DCache.scala 36:26]
  reg  way0Age_24; // @[DCache.scala 36:26]
  reg  way0Age_25; // @[DCache.scala 36:26]
  reg  way0Age_26; // @[DCache.scala 36:26]
  reg  way0Age_27; // @[DCache.scala 36:26]
  reg  way0Age_28; // @[DCache.scala 36:26]
  reg  way0Age_29; // @[DCache.scala 36:26]
  reg  way0Age_30; // @[DCache.scala 36:26]
  reg  way0Age_31; // @[DCache.scala 36:26]
  reg  way0Age_32; // @[DCache.scala 36:26]
  reg  way0Age_33; // @[DCache.scala 36:26]
  reg  way0Age_34; // @[DCache.scala 36:26]
  reg  way0Age_35; // @[DCache.scala 36:26]
  reg  way0Age_36; // @[DCache.scala 36:26]
  reg  way0Age_37; // @[DCache.scala 36:26]
  reg  way0Age_38; // @[DCache.scala 36:26]
  reg  way0Age_39; // @[DCache.scala 36:26]
  reg  way0Age_40; // @[DCache.scala 36:26]
  reg  way0Age_41; // @[DCache.scala 36:26]
  reg  way0Age_42; // @[DCache.scala 36:26]
  reg  way0Age_43; // @[DCache.scala 36:26]
  reg  way0Age_44; // @[DCache.scala 36:26]
  reg  way0Age_45; // @[DCache.scala 36:26]
  reg  way0Age_46; // @[DCache.scala 36:26]
  reg  way0Age_47; // @[DCache.scala 36:26]
  reg  way0Age_48; // @[DCache.scala 36:26]
  reg  way0Age_49; // @[DCache.scala 36:26]
  reg  way0Age_50; // @[DCache.scala 36:26]
  reg  way0Age_51; // @[DCache.scala 36:26]
  reg  way0Age_52; // @[DCache.scala 36:26]
  reg  way0Age_53; // @[DCache.scala 36:26]
  reg  way0Age_54; // @[DCache.scala 36:26]
  reg  way0Age_55; // @[DCache.scala 36:26]
  reg  way0Age_56; // @[DCache.scala 36:26]
  reg  way0Age_57; // @[DCache.scala 36:26]
  reg  way0Age_58; // @[DCache.scala 36:26]
  reg  way0Age_59; // @[DCache.scala 36:26]
  reg  way0Age_60; // @[DCache.scala 36:26]
  reg  way0Age_61; // @[DCache.scala 36:26]
  reg  way0Age_62; // @[DCache.scala 36:26]
  reg  way0Age_63; // @[DCache.scala 36:26]
  reg  way0Age_64; // @[DCache.scala 36:26]
  reg  way0Age_65; // @[DCache.scala 36:26]
  reg  way0Age_66; // @[DCache.scala 36:26]
  reg  way0Age_67; // @[DCache.scala 36:26]
  reg  way0Age_68; // @[DCache.scala 36:26]
  reg  way0Age_69; // @[DCache.scala 36:26]
  reg  way0Age_70; // @[DCache.scala 36:26]
  reg  way0Age_71; // @[DCache.scala 36:26]
  reg  way0Age_72; // @[DCache.scala 36:26]
  reg  way0Age_73; // @[DCache.scala 36:26]
  reg  way0Age_74; // @[DCache.scala 36:26]
  reg  way0Age_75; // @[DCache.scala 36:26]
  reg  way0Age_76; // @[DCache.scala 36:26]
  reg  way0Age_77; // @[DCache.scala 36:26]
  reg  way0Age_78; // @[DCache.scala 36:26]
  reg  way0Age_79; // @[DCache.scala 36:26]
  reg  way0Age_80; // @[DCache.scala 36:26]
  reg  way0Age_81; // @[DCache.scala 36:26]
  reg  way0Age_82; // @[DCache.scala 36:26]
  reg  way0Age_83; // @[DCache.scala 36:26]
  reg  way0Age_84; // @[DCache.scala 36:26]
  reg  way0Age_85; // @[DCache.scala 36:26]
  reg  way0Age_86; // @[DCache.scala 36:26]
  reg  way0Age_87; // @[DCache.scala 36:26]
  reg  way0Age_88; // @[DCache.scala 36:26]
  reg  way0Age_89; // @[DCache.scala 36:26]
  reg  way0Age_90; // @[DCache.scala 36:26]
  reg  way0Age_91; // @[DCache.scala 36:26]
  reg  way0Age_92; // @[DCache.scala 36:26]
  reg  way0Age_93; // @[DCache.scala 36:26]
  reg  way0Age_94; // @[DCache.scala 36:26]
  reg  way0Age_95; // @[DCache.scala 36:26]
  reg  way0Age_96; // @[DCache.scala 36:26]
  reg  way0Age_97; // @[DCache.scala 36:26]
  reg  way0Age_98; // @[DCache.scala 36:26]
  reg  way0Age_99; // @[DCache.scala 36:26]
  reg  way0Age_100; // @[DCache.scala 36:26]
  reg  way0Age_101; // @[DCache.scala 36:26]
  reg  way0Age_102; // @[DCache.scala 36:26]
  reg  way0Age_103; // @[DCache.scala 36:26]
  reg  way0Age_104; // @[DCache.scala 36:26]
  reg  way0Age_105; // @[DCache.scala 36:26]
  reg  way0Age_106; // @[DCache.scala 36:26]
  reg  way0Age_107; // @[DCache.scala 36:26]
  reg  way0Age_108; // @[DCache.scala 36:26]
  reg  way0Age_109; // @[DCache.scala 36:26]
  reg  way0Age_110; // @[DCache.scala 36:26]
  reg  way0Age_111; // @[DCache.scala 36:26]
  reg  way0Age_112; // @[DCache.scala 36:26]
  reg  way0Age_113; // @[DCache.scala 36:26]
  reg  way0Age_114; // @[DCache.scala 36:26]
  reg  way0Age_115; // @[DCache.scala 36:26]
  reg  way0Age_116; // @[DCache.scala 36:26]
  reg  way0Age_117; // @[DCache.scala 36:26]
  reg  way0Age_118; // @[DCache.scala 36:26]
  reg  way0Age_119; // @[DCache.scala 36:26]
  reg  way0Age_120; // @[DCache.scala 36:26]
  reg  way0Age_121; // @[DCache.scala 36:26]
  reg  way0Age_122; // @[DCache.scala 36:26]
  reg  way0Age_123; // @[DCache.scala 36:26]
  reg  way0Age_124; // @[DCache.scala 36:26]
  reg  way0Age_125; // @[DCache.scala 36:26]
  reg  way0Age_126; // @[DCache.scala 36:26]
  reg  way0Age_127; // @[DCache.scala 36:26]
  reg  way0Dirty_0; // @[DCache.scala 37:26]
  reg  way0Dirty_1; // @[DCache.scala 37:26]
  reg  way0Dirty_2; // @[DCache.scala 37:26]
  reg  way0Dirty_3; // @[DCache.scala 37:26]
  reg  way0Dirty_4; // @[DCache.scala 37:26]
  reg  way0Dirty_5; // @[DCache.scala 37:26]
  reg  way0Dirty_6; // @[DCache.scala 37:26]
  reg  way0Dirty_7; // @[DCache.scala 37:26]
  reg  way0Dirty_8; // @[DCache.scala 37:26]
  reg  way0Dirty_9; // @[DCache.scala 37:26]
  reg  way0Dirty_10; // @[DCache.scala 37:26]
  reg  way0Dirty_11; // @[DCache.scala 37:26]
  reg  way0Dirty_12; // @[DCache.scala 37:26]
  reg  way0Dirty_13; // @[DCache.scala 37:26]
  reg  way0Dirty_14; // @[DCache.scala 37:26]
  reg  way0Dirty_15; // @[DCache.scala 37:26]
  reg  way0Dirty_16; // @[DCache.scala 37:26]
  reg  way0Dirty_17; // @[DCache.scala 37:26]
  reg  way0Dirty_18; // @[DCache.scala 37:26]
  reg  way0Dirty_19; // @[DCache.scala 37:26]
  reg  way0Dirty_20; // @[DCache.scala 37:26]
  reg  way0Dirty_21; // @[DCache.scala 37:26]
  reg  way0Dirty_22; // @[DCache.scala 37:26]
  reg  way0Dirty_23; // @[DCache.scala 37:26]
  reg  way0Dirty_24; // @[DCache.scala 37:26]
  reg  way0Dirty_25; // @[DCache.scala 37:26]
  reg  way0Dirty_26; // @[DCache.scala 37:26]
  reg  way0Dirty_27; // @[DCache.scala 37:26]
  reg  way0Dirty_28; // @[DCache.scala 37:26]
  reg  way0Dirty_29; // @[DCache.scala 37:26]
  reg  way0Dirty_30; // @[DCache.scala 37:26]
  reg  way0Dirty_31; // @[DCache.scala 37:26]
  reg  way0Dirty_32; // @[DCache.scala 37:26]
  reg  way0Dirty_33; // @[DCache.scala 37:26]
  reg  way0Dirty_34; // @[DCache.scala 37:26]
  reg  way0Dirty_35; // @[DCache.scala 37:26]
  reg  way0Dirty_36; // @[DCache.scala 37:26]
  reg  way0Dirty_37; // @[DCache.scala 37:26]
  reg  way0Dirty_38; // @[DCache.scala 37:26]
  reg  way0Dirty_39; // @[DCache.scala 37:26]
  reg  way0Dirty_40; // @[DCache.scala 37:26]
  reg  way0Dirty_41; // @[DCache.scala 37:26]
  reg  way0Dirty_42; // @[DCache.scala 37:26]
  reg  way0Dirty_43; // @[DCache.scala 37:26]
  reg  way0Dirty_44; // @[DCache.scala 37:26]
  reg  way0Dirty_45; // @[DCache.scala 37:26]
  reg  way0Dirty_46; // @[DCache.scala 37:26]
  reg  way0Dirty_47; // @[DCache.scala 37:26]
  reg  way0Dirty_48; // @[DCache.scala 37:26]
  reg  way0Dirty_49; // @[DCache.scala 37:26]
  reg  way0Dirty_50; // @[DCache.scala 37:26]
  reg  way0Dirty_51; // @[DCache.scala 37:26]
  reg  way0Dirty_52; // @[DCache.scala 37:26]
  reg  way0Dirty_53; // @[DCache.scala 37:26]
  reg  way0Dirty_54; // @[DCache.scala 37:26]
  reg  way0Dirty_55; // @[DCache.scala 37:26]
  reg  way0Dirty_56; // @[DCache.scala 37:26]
  reg  way0Dirty_57; // @[DCache.scala 37:26]
  reg  way0Dirty_58; // @[DCache.scala 37:26]
  reg  way0Dirty_59; // @[DCache.scala 37:26]
  reg  way0Dirty_60; // @[DCache.scala 37:26]
  reg  way0Dirty_61; // @[DCache.scala 37:26]
  reg  way0Dirty_62; // @[DCache.scala 37:26]
  reg  way0Dirty_63; // @[DCache.scala 37:26]
  reg  way0Dirty_64; // @[DCache.scala 37:26]
  reg  way0Dirty_65; // @[DCache.scala 37:26]
  reg  way0Dirty_66; // @[DCache.scala 37:26]
  reg  way0Dirty_67; // @[DCache.scala 37:26]
  reg  way0Dirty_68; // @[DCache.scala 37:26]
  reg  way0Dirty_69; // @[DCache.scala 37:26]
  reg  way0Dirty_70; // @[DCache.scala 37:26]
  reg  way0Dirty_71; // @[DCache.scala 37:26]
  reg  way0Dirty_72; // @[DCache.scala 37:26]
  reg  way0Dirty_73; // @[DCache.scala 37:26]
  reg  way0Dirty_74; // @[DCache.scala 37:26]
  reg  way0Dirty_75; // @[DCache.scala 37:26]
  reg  way0Dirty_76; // @[DCache.scala 37:26]
  reg  way0Dirty_77; // @[DCache.scala 37:26]
  reg  way0Dirty_78; // @[DCache.scala 37:26]
  reg  way0Dirty_79; // @[DCache.scala 37:26]
  reg  way0Dirty_80; // @[DCache.scala 37:26]
  reg  way0Dirty_81; // @[DCache.scala 37:26]
  reg  way0Dirty_82; // @[DCache.scala 37:26]
  reg  way0Dirty_83; // @[DCache.scala 37:26]
  reg  way0Dirty_84; // @[DCache.scala 37:26]
  reg  way0Dirty_85; // @[DCache.scala 37:26]
  reg  way0Dirty_86; // @[DCache.scala 37:26]
  reg  way0Dirty_87; // @[DCache.scala 37:26]
  reg  way0Dirty_88; // @[DCache.scala 37:26]
  reg  way0Dirty_89; // @[DCache.scala 37:26]
  reg  way0Dirty_90; // @[DCache.scala 37:26]
  reg  way0Dirty_91; // @[DCache.scala 37:26]
  reg  way0Dirty_92; // @[DCache.scala 37:26]
  reg  way0Dirty_93; // @[DCache.scala 37:26]
  reg  way0Dirty_94; // @[DCache.scala 37:26]
  reg  way0Dirty_95; // @[DCache.scala 37:26]
  reg  way0Dirty_96; // @[DCache.scala 37:26]
  reg  way0Dirty_97; // @[DCache.scala 37:26]
  reg  way0Dirty_98; // @[DCache.scala 37:26]
  reg  way0Dirty_99; // @[DCache.scala 37:26]
  reg  way0Dirty_100; // @[DCache.scala 37:26]
  reg  way0Dirty_101; // @[DCache.scala 37:26]
  reg  way0Dirty_102; // @[DCache.scala 37:26]
  reg  way0Dirty_103; // @[DCache.scala 37:26]
  reg  way0Dirty_104; // @[DCache.scala 37:26]
  reg  way0Dirty_105; // @[DCache.scala 37:26]
  reg  way0Dirty_106; // @[DCache.scala 37:26]
  reg  way0Dirty_107; // @[DCache.scala 37:26]
  reg  way0Dirty_108; // @[DCache.scala 37:26]
  reg  way0Dirty_109; // @[DCache.scala 37:26]
  reg  way0Dirty_110; // @[DCache.scala 37:26]
  reg  way0Dirty_111; // @[DCache.scala 37:26]
  reg  way0Dirty_112; // @[DCache.scala 37:26]
  reg  way0Dirty_113; // @[DCache.scala 37:26]
  reg  way0Dirty_114; // @[DCache.scala 37:26]
  reg  way0Dirty_115; // @[DCache.scala 37:26]
  reg  way0Dirty_116; // @[DCache.scala 37:26]
  reg  way0Dirty_117; // @[DCache.scala 37:26]
  reg  way0Dirty_118; // @[DCache.scala 37:26]
  reg  way0Dirty_119; // @[DCache.scala 37:26]
  reg  way0Dirty_120; // @[DCache.scala 37:26]
  reg  way0Dirty_121; // @[DCache.scala 37:26]
  reg  way0Dirty_122; // @[DCache.scala 37:26]
  reg  way0Dirty_123; // @[DCache.scala 37:26]
  reg  way0Dirty_124; // @[DCache.scala 37:26]
  reg  way0Dirty_125; // @[DCache.scala 37:26]
  reg  way0Dirty_126; // @[DCache.scala 37:26]
  reg  way0Dirty_127; // @[DCache.scala 37:26]
  reg  way1V_0; // @[DCache.scala 39:26]
  reg  way1V_1; // @[DCache.scala 39:26]
  reg  way1V_2; // @[DCache.scala 39:26]
  reg  way1V_3; // @[DCache.scala 39:26]
  reg  way1V_4; // @[DCache.scala 39:26]
  reg  way1V_5; // @[DCache.scala 39:26]
  reg  way1V_6; // @[DCache.scala 39:26]
  reg  way1V_7; // @[DCache.scala 39:26]
  reg  way1V_8; // @[DCache.scala 39:26]
  reg  way1V_9; // @[DCache.scala 39:26]
  reg  way1V_10; // @[DCache.scala 39:26]
  reg  way1V_11; // @[DCache.scala 39:26]
  reg  way1V_12; // @[DCache.scala 39:26]
  reg  way1V_13; // @[DCache.scala 39:26]
  reg  way1V_14; // @[DCache.scala 39:26]
  reg  way1V_15; // @[DCache.scala 39:26]
  reg  way1V_16; // @[DCache.scala 39:26]
  reg  way1V_17; // @[DCache.scala 39:26]
  reg  way1V_18; // @[DCache.scala 39:26]
  reg  way1V_19; // @[DCache.scala 39:26]
  reg  way1V_20; // @[DCache.scala 39:26]
  reg  way1V_21; // @[DCache.scala 39:26]
  reg  way1V_22; // @[DCache.scala 39:26]
  reg  way1V_23; // @[DCache.scala 39:26]
  reg  way1V_24; // @[DCache.scala 39:26]
  reg  way1V_25; // @[DCache.scala 39:26]
  reg  way1V_26; // @[DCache.scala 39:26]
  reg  way1V_27; // @[DCache.scala 39:26]
  reg  way1V_28; // @[DCache.scala 39:26]
  reg  way1V_29; // @[DCache.scala 39:26]
  reg  way1V_30; // @[DCache.scala 39:26]
  reg  way1V_31; // @[DCache.scala 39:26]
  reg  way1V_32; // @[DCache.scala 39:26]
  reg  way1V_33; // @[DCache.scala 39:26]
  reg  way1V_34; // @[DCache.scala 39:26]
  reg  way1V_35; // @[DCache.scala 39:26]
  reg  way1V_36; // @[DCache.scala 39:26]
  reg  way1V_37; // @[DCache.scala 39:26]
  reg  way1V_38; // @[DCache.scala 39:26]
  reg  way1V_39; // @[DCache.scala 39:26]
  reg  way1V_40; // @[DCache.scala 39:26]
  reg  way1V_41; // @[DCache.scala 39:26]
  reg  way1V_42; // @[DCache.scala 39:26]
  reg  way1V_43; // @[DCache.scala 39:26]
  reg  way1V_44; // @[DCache.scala 39:26]
  reg  way1V_45; // @[DCache.scala 39:26]
  reg  way1V_46; // @[DCache.scala 39:26]
  reg  way1V_47; // @[DCache.scala 39:26]
  reg  way1V_48; // @[DCache.scala 39:26]
  reg  way1V_49; // @[DCache.scala 39:26]
  reg  way1V_50; // @[DCache.scala 39:26]
  reg  way1V_51; // @[DCache.scala 39:26]
  reg  way1V_52; // @[DCache.scala 39:26]
  reg  way1V_53; // @[DCache.scala 39:26]
  reg  way1V_54; // @[DCache.scala 39:26]
  reg  way1V_55; // @[DCache.scala 39:26]
  reg  way1V_56; // @[DCache.scala 39:26]
  reg  way1V_57; // @[DCache.scala 39:26]
  reg  way1V_58; // @[DCache.scala 39:26]
  reg  way1V_59; // @[DCache.scala 39:26]
  reg  way1V_60; // @[DCache.scala 39:26]
  reg  way1V_61; // @[DCache.scala 39:26]
  reg  way1V_62; // @[DCache.scala 39:26]
  reg  way1V_63; // @[DCache.scala 39:26]
  reg  way1V_64; // @[DCache.scala 39:26]
  reg  way1V_65; // @[DCache.scala 39:26]
  reg  way1V_66; // @[DCache.scala 39:26]
  reg  way1V_67; // @[DCache.scala 39:26]
  reg  way1V_68; // @[DCache.scala 39:26]
  reg  way1V_69; // @[DCache.scala 39:26]
  reg  way1V_70; // @[DCache.scala 39:26]
  reg  way1V_71; // @[DCache.scala 39:26]
  reg  way1V_72; // @[DCache.scala 39:26]
  reg  way1V_73; // @[DCache.scala 39:26]
  reg  way1V_74; // @[DCache.scala 39:26]
  reg  way1V_75; // @[DCache.scala 39:26]
  reg  way1V_76; // @[DCache.scala 39:26]
  reg  way1V_77; // @[DCache.scala 39:26]
  reg  way1V_78; // @[DCache.scala 39:26]
  reg  way1V_79; // @[DCache.scala 39:26]
  reg  way1V_80; // @[DCache.scala 39:26]
  reg  way1V_81; // @[DCache.scala 39:26]
  reg  way1V_82; // @[DCache.scala 39:26]
  reg  way1V_83; // @[DCache.scala 39:26]
  reg  way1V_84; // @[DCache.scala 39:26]
  reg  way1V_85; // @[DCache.scala 39:26]
  reg  way1V_86; // @[DCache.scala 39:26]
  reg  way1V_87; // @[DCache.scala 39:26]
  reg  way1V_88; // @[DCache.scala 39:26]
  reg  way1V_89; // @[DCache.scala 39:26]
  reg  way1V_90; // @[DCache.scala 39:26]
  reg  way1V_91; // @[DCache.scala 39:26]
  reg  way1V_92; // @[DCache.scala 39:26]
  reg  way1V_93; // @[DCache.scala 39:26]
  reg  way1V_94; // @[DCache.scala 39:26]
  reg  way1V_95; // @[DCache.scala 39:26]
  reg  way1V_96; // @[DCache.scala 39:26]
  reg  way1V_97; // @[DCache.scala 39:26]
  reg  way1V_98; // @[DCache.scala 39:26]
  reg  way1V_99; // @[DCache.scala 39:26]
  reg  way1V_100; // @[DCache.scala 39:26]
  reg  way1V_101; // @[DCache.scala 39:26]
  reg  way1V_102; // @[DCache.scala 39:26]
  reg  way1V_103; // @[DCache.scala 39:26]
  reg  way1V_104; // @[DCache.scala 39:26]
  reg  way1V_105; // @[DCache.scala 39:26]
  reg  way1V_106; // @[DCache.scala 39:26]
  reg  way1V_107; // @[DCache.scala 39:26]
  reg  way1V_108; // @[DCache.scala 39:26]
  reg  way1V_109; // @[DCache.scala 39:26]
  reg  way1V_110; // @[DCache.scala 39:26]
  reg  way1V_111; // @[DCache.scala 39:26]
  reg  way1V_112; // @[DCache.scala 39:26]
  reg  way1V_113; // @[DCache.scala 39:26]
  reg  way1V_114; // @[DCache.scala 39:26]
  reg  way1V_115; // @[DCache.scala 39:26]
  reg  way1V_116; // @[DCache.scala 39:26]
  reg  way1V_117; // @[DCache.scala 39:26]
  reg  way1V_118; // @[DCache.scala 39:26]
  reg  way1V_119; // @[DCache.scala 39:26]
  reg  way1V_120; // @[DCache.scala 39:26]
  reg  way1V_121; // @[DCache.scala 39:26]
  reg  way1V_122; // @[DCache.scala 39:26]
  reg  way1V_123; // @[DCache.scala 39:26]
  reg  way1V_124; // @[DCache.scala 39:26]
  reg  way1V_125; // @[DCache.scala 39:26]
  reg  way1V_126; // @[DCache.scala 39:26]
  reg  way1V_127; // @[DCache.scala 39:26]
  reg [20:0] way1Tag_0; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_1; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_2; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_3; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_4; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_5; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_6; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_7; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_8; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_9; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_10; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_11; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_12; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_13; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_14; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_15; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_16; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_17; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_18; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_19; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_20; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_21; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_22; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_23; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_24; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_25; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_26; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_27; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_28; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_29; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_30; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_31; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_32; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_33; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_34; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_35; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_36; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_37; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_38; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_39; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_40; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_41; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_42; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_43; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_44; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_45; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_46; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_47; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_48; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_49; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_50; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_51; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_52; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_53; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_54; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_55; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_56; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_57; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_58; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_59; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_60; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_61; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_62; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_63; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_64; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_65; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_66; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_67; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_68; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_69; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_70; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_71; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_72; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_73; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_74; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_75; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_76; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_77; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_78; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_79; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_80; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_81; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_82; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_83; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_84; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_85; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_86; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_87; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_88; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_89; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_90; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_91; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_92; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_93; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_94; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_95; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_96; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_97; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_98; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_99; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_100; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_101; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_102; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_103; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_104; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_105; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_106; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_107; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_108; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_109; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_110; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_111; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_112; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_113; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_114; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_115; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_116; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_117; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_118; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_119; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_120; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_121; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_122; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_123; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_124; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_125; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_126; // @[DCache.scala 40:26]
  reg [20:0] way1Tag_127; // @[DCache.scala 40:26]
  reg  way1Age_0; // @[DCache.scala 42:26]
  reg  way1Age_1; // @[DCache.scala 42:26]
  reg  way1Age_2; // @[DCache.scala 42:26]
  reg  way1Age_3; // @[DCache.scala 42:26]
  reg  way1Age_4; // @[DCache.scala 42:26]
  reg  way1Age_5; // @[DCache.scala 42:26]
  reg  way1Age_6; // @[DCache.scala 42:26]
  reg  way1Age_7; // @[DCache.scala 42:26]
  reg  way1Age_8; // @[DCache.scala 42:26]
  reg  way1Age_9; // @[DCache.scala 42:26]
  reg  way1Age_10; // @[DCache.scala 42:26]
  reg  way1Age_11; // @[DCache.scala 42:26]
  reg  way1Age_12; // @[DCache.scala 42:26]
  reg  way1Age_13; // @[DCache.scala 42:26]
  reg  way1Age_14; // @[DCache.scala 42:26]
  reg  way1Age_15; // @[DCache.scala 42:26]
  reg  way1Age_16; // @[DCache.scala 42:26]
  reg  way1Age_17; // @[DCache.scala 42:26]
  reg  way1Age_18; // @[DCache.scala 42:26]
  reg  way1Age_19; // @[DCache.scala 42:26]
  reg  way1Age_20; // @[DCache.scala 42:26]
  reg  way1Age_21; // @[DCache.scala 42:26]
  reg  way1Age_22; // @[DCache.scala 42:26]
  reg  way1Age_23; // @[DCache.scala 42:26]
  reg  way1Age_24; // @[DCache.scala 42:26]
  reg  way1Age_25; // @[DCache.scala 42:26]
  reg  way1Age_26; // @[DCache.scala 42:26]
  reg  way1Age_27; // @[DCache.scala 42:26]
  reg  way1Age_28; // @[DCache.scala 42:26]
  reg  way1Age_29; // @[DCache.scala 42:26]
  reg  way1Age_30; // @[DCache.scala 42:26]
  reg  way1Age_31; // @[DCache.scala 42:26]
  reg  way1Age_32; // @[DCache.scala 42:26]
  reg  way1Age_33; // @[DCache.scala 42:26]
  reg  way1Age_34; // @[DCache.scala 42:26]
  reg  way1Age_35; // @[DCache.scala 42:26]
  reg  way1Age_36; // @[DCache.scala 42:26]
  reg  way1Age_37; // @[DCache.scala 42:26]
  reg  way1Age_38; // @[DCache.scala 42:26]
  reg  way1Age_39; // @[DCache.scala 42:26]
  reg  way1Age_40; // @[DCache.scala 42:26]
  reg  way1Age_41; // @[DCache.scala 42:26]
  reg  way1Age_42; // @[DCache.scala 42:26]
  reg  way1Age_43; // @[DCache.scala 42:26]
  reg  way1Age_44; // @[DCache.scala 42:26]
  reg  way1Age_45; // @[DCache.scala 42:26]
  reg  way1Age_46; // @[DCache.scala 42:26]
  reg  way1Age_47; // @[DCache.scala 42:26]
  reg  way1Age_48; // @[DCache.scala 42:26]
  reg  way1Age_49; // @[DCache.scala 42:26]
  reg  way1Age_50; // @[DCache.scala 42:26]
  reg  way1Age_51; // @[DCache.scala 42:26]
  reg  way1Age_52; // @[DCache.scala 42:26]
  reg  way1Age_53; // @[DCache.scala 42:26]
  reg  way1Age_54; // @[DCache.scala 42:26]
  reg  way1Age_55; // @[DCache.scala 42:26]
  reg  way1Age_56; // @[DCache.scala 42:26]
  reg  way1Age_57; // @[DCache.scala 42:26]
  reg  way1Age_58; // @[DCache.scala 42:26]
  reg  way1Age_59; // @[DCache.scala 42:26]
  reg  way1Age_60; // @[DCache.scala 42:26]
  reg  way1Age_61; // @[DCache.scala 42:26]
  reg  way1Age_62; // @[DCache.scala 42:26]
  reg  way1Age_63; // @[DCache.scala 42:26]
  reg  way1Age_64; // @[DCache.scala 42:26]
  reg  way1Age_65; // @[DCache.scala 42:26]
  reg  way1Age_66; // @[DCache.scala 42:26]
  reg  way1Age_67; // @[DCache.scala 42:26]
  reg  way1Age_68; // @[DCache.scala 42:26]
  reg  way1Age_69; // @[DCache.scala 42:26]
  reg  way1Age_70; // @[DCache.scala 42:26]
  reg  way1Age_71; // @[DCache.scala 42:26]
  reg  way1Age_72; // @[DCache.scala 42:26]
  reg  way1Age_73; // @[DCache.scala 42:26]
  reg  way1Age_74; // @[DCache.scala 42:26]
  reg  way1Age_75; // @[DCache.scala 42:26]
  reg  way1Age_76; // @[DCache.scala 42:26]
  reg  way1Age_77; // @[DCache.scala 42:26]
  reg  way1Age_78; // @[DCache.scala 42:26]
  reg  way1Age_79; // @[DCache.scala 42:26]
  reg  way1Age_80; // @[DCache.scala 42:26]
  reg  way1Age_81; // @[DCache.scala 42:26]
  reg  way1Age_82; // @[DCache.scala 42:26]
  reg  way1Age_83; // @[DCache.scala 42:26]
  reg  way1Age_84; // @[DCache.scala 42:26]
  reg  way1Age_85; // @[DCache.scala 42:26]
  reg  way1Age_86; // @[DCache.scala 42:26]
  reg  way1Age_87; // @[DCache.scala 42:26]
  reg  way1Age_88; // @[DCache.scala 42:26]
  reg  way1Age_89; // @[DCache.scala 42:26]
  reg  way1Age_90; // @[DCache.scala 42:26]
  reg  way1Age_91; // @[DCache.scala 42:26]
  reg  way1Age_92; // @[DCache.scala 42:26]
  reg  way1Age_93; // @[DCache.scala 42:26]
  reg  way1Age_94; // @[DCache.scala 42:26]
  reg  way1Age_95; // @[DCache.scala 42:26]
  reg  way1Age_96; // @[DCache.scala 42:26]
  reg  way1Age_97; // @[DCache.scala 42:26]
  reg  way1Age_98; // @[DCache.scala 42:26]
  reg  way1Age_99; // @[DCache.scala 42:26]
  reg  way1Age_100; // @[DCache.scala 42:26]
  reg  way1Age_101; // @[DCache.scala 42:26]
  reg  way1Age_102; // @[DCache.scala 42:26]
  reg  way1Age_103; // @[DCache.scala 42:26]
  reg  way1Age_104; // @[DCache.scala 42:26]
  reg  way1Age_105; // @[DCache.scala 42:26]
  reg  way1Age_106; // @[DCache.scala 42:26]
  reg  way1Age_107; // @[DCache.scala 42:26]
  reg  way1Age_108; // @[DCache.scala 42:26]
  reg  way1Age_109; // @[DCache.scala 42:26]
  reg  way1Age_110; // @[DCache.scala 42:26]
  reg  way1Age_111; // @[DCache.scala 42:26]
  reg  way1Age_112; // @[DCache.scala 42:26]
  reg  way1Age_113; // @[DCache.scala 42:26]
  reg  way1Age_114; // @[DCache.scala 42:26]
  reg  way1Age_115; // @[DCache.scala 42:26]
  reg  way1Age_116; // @[DCache.scala 42:26]
  reg  way1Age_117; // @[DCache.scala 42:26]
  reg  way1Age_118; // @[DCache.scala 42:26]
  reg  way1Age_119; // @[DCache.scala 42:26]
  reg  way1Age_120; // @[DCache.scala 42:26]
  reg  way1Age_121; // @[DCache.scala 42:26]
  reg  way1Age_122; // @[DCache.scala 42:26]
  reg  way1Age_123; // @[DCache.scala 42:26]
  reg  way1Age_124; // @[DCache.scala 42:26]
  reg  way1Age_125; // @[DCache.scala 42:26]
  reg  way1Age_126; // @[DCache.scala 42:26]
  reg  way1Age_127; // @[DCache.scala 42:26]
  reg  way1Dirty_0; // @[DCache.scala 43:26]
  reg  way1Dirty_1; // @[DCache.scala 43:26]
  reg  way1Dirty_2; // @[DCache.scala 43:26]
  reg  way1Dirty_3; // @[DCache.scala 43:26]
  reg  way1Dirty_4; // @[DCache.scala 43:26]
  reg  way1Dirty_5; // @[DCache.scala 43:26]
  reg  way1Dirty_6; // @[DCache.scala 43:26]
  reg  way1Dirty_7; // @[DCache.scala 43:26]
  reg  way1Dirty_8; // @[DCache.scala 43:26]
  reg  way1Dirty_9; // @[DCache.scala 43:26]
  reg  way1Dirty_10; // @[DCache.scala 43:26]
  reg  way1Dirty_11; // @[DCache.scala 43:26]
  reg  way1Dirty_12; // @[DCache.scala 43:26]
  reg  way1Dirty_13; // @[DCache.scala 43:26]
  reg  way1Dirty_14; // @[DCache.scala 43:26]
  reg  way1Dirty_15; // @[DCache.scala 43:26]
  reg  way1Dirty_16; // @[DCache.scala 43:26]
  reg  way1Dirty_17; // @[DCache.scala 43:26]
  reg  way1Dirty_18; // @[DCache.scala 43:26]
  reg  way1Dirty_19; // @[DCache.scala 43:26]
  reg  way1Dirty_20; // @[DCache.scala 43:26]
  reg  way1Dirty_21; // @[DCache.scala 43:26]
  reg  way1Dirty_22; // @[DCache.scala 43:26]
  reg  way1Dirty_23; // @[DCache.scala 43:26]
  reg  way1Dirty_24; // @[DCache.scala 43:26]
  reg  way1Dirty_25; // @[DCache.scala 43:26]
  reg  way1Dirty_26; // @[DCache.scala 43:26]
  reg  way1Dirty_27; // @[DCache.scala 43:26]
  reg  way1Dirty_28; // @[DCache.scala 43:26]
  reg  way1Dirty_29; // @[DCache.scala 43:26]
  reg  way1Dirty_30; // @[DCache.scala 43:26]
  reg  way1Dirty_31; // @[DCache.scala 43:26]
  reg  way1Dirty_32; // @[DCache.scala 43:26]
  reg  way1Dirty_33; // @[DCache.scala 43:26]
  reg  way1Dirty_34; // @[DCache.scala 43:26]
  reg  way1Dirty_35; // @[DCache.scala 43:26]
  reg  way1Dirty_36; // @[DCache.scala 43:26]
  reg  way1Dirty_37; // @[DCache.scala 43:26]
  reg  way1Dirty_38; // @[DCache.scala 43:26]
  reg  way1Dirty_39; // @[DCache.scala 43:26]
  reg  way1Dirty_40; // @[DCache.scala 43:26]
  reg  way1Dirty_41; // @[DCache.scala 43:26]
  reg  way1Dirty_42; // @[DCache.scala 43:26]
  reg  way1Dirty_43; // @[DCache.scala 43:26]
  reg  way1Dirty_44; // @[DCache.scala 43:26]
  reg  way1Dirty_45; // @[DCache.scala 43:26]
  reg  way1Dirty_46; // @[DCache.scala 43:26]
  reg  way1Dirty_47; // @[DCache.scala 43:26]
  reg  way1Dirty_48; // @[DCache.scala 43:26]
  reg  way1Dirty_49; // @[DCache.scala 43:26]
  reg  way1Dirty_50; // @[DCache.scala 43:26]
  reg  way1Dirty_51; // @[DCache.scala 43:26]
  reg  way1Dirty_52; // @[DCache.scala 43:26]
  reg  way1Dirty_53; // @[DCache.scala 43:26]
  reg  way1Dirty_54; // @[DCache.scala 43:26]
  reg  way1Dirty_55; // @[DCache.scala 43:26]
  reg  way1Dirty_56; // @[DCache.scala 43:26]
  reg  way1Dirty_57; // @[DCache.scala 43:26]
  reg  way1Dirty_58; // @[DCache.scala 43:26]
  reg  way1Dirty_59; // @[DCache.scala 43:26]
  reg  way1Dirty_60; // @[DCache.scala 43:26]
  reg  way1Dirty_61; // @[DCache.scala 43:26]
  reg  way1Dirty_62; // @[DCache.scala 43:26]
  reg  way1Dirty_63; // @[DCache.scala 43:26]
  reg  way1Dirty_64; // @[DCache.scala 43:26]
  reg  way1Dirty_65; // @[DCache.scala 43:26]
  reg  way1Dirty_66; // @[DCache.scala 43:26]
  reg  way1Dirty_67; // @[DCache.scala 43:26]
  reg  way1Dirty_68; // @[DCache.scala 43:26]
  reg  way1Dirty_69; // @[DCache.scala 43:26]
  reg  way1Dirty_70; // @[DCache.scala 43:26]
  reg  way1Dirty_71; // @[DCache.scala 43:26]
  reg  way1Dirty_72; // @[DCache.scala 43:26]
  reg  way1Dirty_73; // @[DCache.scala 43:26]
  reg  way1Dirty_74; // @[DCache.scala 43:26]
  reg  way1Dirty_75; // @[DCache.scala 43:26]
  reg  way1Dirty_76; // @[DCache.scala 43:26]
  reg  way1Dirty_77; // @[DCache.scala 43:26]
  reg  way1Dirty_78; // @[DCache.scala 43:26]
  reg  way1Dirty_79; // @[DCache.scala 43:26]
  reg  way1Dirty_80; // @[DCache.scala 43:26]
  reg  way1Dirty_81; // @[DCache.scala 43:26]
  reg  way1Dirty_82; // @[DCache.scala 43:26]
  reg  way1Dirty_83; // @[DCache.scala 43:26]
  reg  way1Dirty_84; // @[DCache.scala 43:26]
  reg  way1Dirty_85; // @[DCache.scala 43:26]
  reg  way1Dirty_86; // @[DCache.scala 43:26]
  reg  way1Dirty_87; // @[DCache.scala 43:26]
  reg  way1Dirty_88; // @[DCache.scala 43:26]
  reg  way1Dirty_89; // @[DCache.scala 43:26]
  reg  way1Dirty_90; // @[DCache.scala 43:26]
  reg  way1Dirty_91; // @[DCache.scala 43:26]
  reg  way1Dirty_92; // @[DCache.scala 43:26]
  reg  way1Dirty_93; // @[DCache.scala 43:26]
  reg  way1Dirty_94; // @[DCache.scala 43:26]
  reg  way1Dirty_95; // @[DCache.scala 43:26]
  reg  way1Dirty_96; // @[DCache.scala 43:26]
  reg  way1Dirty_97; // @[DCache.scala 43:26]
  reg  way1Dirty_98; // @[DCache.scala 43:26]
  reg  way1Dirty_99; // @[DCache.scala 43:26]
  reg  way1Dirty_100; // @[DCache.scala 43:26]
  reg  way1Dirty_101; // @[DCache.scala 43:26]
  reg  way1Dirty_102; // @[DCache.scala 43:26]
  reg  way1Dirty_103; // @[DCache.scala 43:26]
  reg  way1Dirty_104; // @[DCache.scala 43:26]
  reg  way1Dirty_105; // @[DCache.scala 43:26]
  reg  way1Dirty_106; // @[DCache.scala 43:26]
  reg  way1Dirty_107; // @[DCache.scala 43:26]
  reg  way1Dirty_108; // @[DCache.scala 43:26]
  reg  way1Dirty_109; // @[DCache.scala 43:26]
  reg  way1Dirty_110; // @[DCache.scala 43:26]
  reg  way1Dirty_111; // @[DCache.scala 43:26]
  reg  way1Dirty_112; // @[DCache.scala 43:26]
  reg  way1Dirty_113; // @[DCache.scala 43:26]
  reg  way1Dirty_114; // @[DCache.scala 43:26]
  reg  way1Dirty_115; // @[DCache.scala 43:26]
  reg  way1Dirty_116; // @[DCache.scala 43:26]
  reg  way1Dirty_117; // @[DCache.scala 43:26]
  reg  way1Dirty_118; // @[DCache.scala 43:26]
  reg  way1Dirty_119; // @[DCache.scala 43:26]
  reg  way1Dirty_120; // @[DCache.scala 43:26]
  reg  way1Dirty_121; // @[DCache.scala 43:26]
  reg  way1Dirty_122; // @[DCache.scala 43:26]
  reg  way1Dirty_123; // @[DCache.scala 43:26]
  reg  way1Dirty_124; // @[DCache.scala 43:26]
  reg  way1Dirty_125; // @[DCache.scala 43:26]
  reg  way1Dirty_126; // @[DCache.scala 43:26]
  reg  way1Dirty_127; // @[DCache.scala 43:26]
  reg [2:0] state; // @[DCache.scala 46:22]
  wire [20:0] reqTag = io_dmem_data_addr[31:11]; // @[DCache.scala 50:27]
  wire [6:0] reqIndex = io_dmem_data_addr[10:4]; // @[DCache.scala 51:27]
  wire [3:0] reqOff = io_dmem_data_addr[3:0]; // @[DCache.scala 52:27]
  wire [7:0] _strbT_T_1 = 8'h1 == io_dmem_data_strb ? 8'hff : 8'h0; // @[Mux.scala 81:58]
  wire [15:0] _strbT_T_3 = 8'h2 == io_dmem_data_strb ? 16'hff00 : {{8'd0}, _strbT_T_1}; // @[Mux.scala 81:58]
  wire [23:0] _strbT_T_5 = 8'h4 == io_dmem_data_strb ? 24'hff0000 : {{8'd0}, _strbT_T_3}; // @[Mux.scala 81:58]
  wire [31:0] _strbT_T_7 = 8'h8 == io_dmem_data_strb ? 32'hff000000 : {{8'd0}, _strbT_T_5}; // @[Mux.scala 81:58]
  wire [39:0] _strbT_T_9 = 8'h10 == io_dmem_data_strb ? 40'hff00000000 : {{8'd0}, _strbT_T_7}; // @[Mux.scala 81:58]
  wire [47:0] _strbT_T_11 = 8'h20 == io_dmem_data_strb ? 48'hff0000000000 : {{8'd0}, _strbT_T_9}; // @[Mux.scala 81:58]
  wire [55:0] _strbT_T_13 = 8'h40 == io_dmem_data_strb ? 56'hff000000000000 : {{8'd0}, _strbT_T_11}; // @[Mux.scala 81:58]
  wire [63:0] _strbT_T_15 = 8'h80 == io_dmem_data_strb ? 64'hff00000000000000 : {{8'd0}, _strbT_T_13}; // @[Mux.scala 81:58]
  wire [63:0] _strbT_T_17 = 8'h3 == io_dmem_data_strb ? 64'hffff : _strbT_T_15; // @[Mux.scala 81:58]
  wire [63:0] _strbT_T_19 = 8'hc == io_dmem_data_strb ? 64'hffff0000 : _strbT_T_17; // @[Mux.scala 81:58]
  wire [63:0] _strbT_T_21 = 8'h30 == io_dmem_data_strb ? 64'hffff00000000 : _strbT_T_19; // @[Mux.scala 81:58]
  wire [63:0] _strbT_T_23 = 8'hc0 == io_dmem_data_strb ? 64'hffff000000000000 : _strbT_T_21; // @[Mux.scala 81:58]
  wire [63:0] _strbT_T_25 = 8'hf == io_dmem_data_strb ? 64'hffffffff : _strbT_T_23; // @[Mux.scala 81:58]
  wire [63:0] _strbT_T_27 = 8'hf0 == io_dmem_data_strb ? 64'hffffffff00000000 : _strbT_T_25; // @[Mux.scala 81:58]
  wire [63:0] strbT = 8'hff == io_dmem_data_strb ? 64'hffffffffffffffff : _strbT_T_27; // @[Mux.scala 81:58]
  wire [127:0] _valid_strb_T_1 = {strbT,64'h0}; // @[Cat.scala 31:58]
  wire [127:0] _valid_strb_T_2 = {64'h0,strbT}; // @[Cat.scala 31:58]
  wire [127:0] valid_strb = reqOff[3] ? _valid_strb_T_1 : _valid_strb_T_2; // @[DCache.scala 72:24]
  wire [2:0] _GEN_1 = ~io_dmem_data_req ? 3'h6 : 3'h5; // @[DCache.scala 85:40 86:17 88:17]
  wire  _GEN_142 = 7'h1 == reqIndex ? way0V_1 : way0V_0; // @[DCache.scala 124:{33,33}]
  wire  _GEN_143 = 7'h2 == reqIndex ? way0V_2 : _GEN_142; // @[DCache.scala 124:{33,33}]
  wire  _GEN_144 = 7'h3 == reqIndex ? way0V_3 : _GEN_143; // @[DCache.scala 124:{33,33}]
  wire  _GEN_145 = 7'h4 == reqIndex ? way0V_4 : _GEN_144; // @[DCache.scala 124:{33,33}]
  wire  _GEN_146 = 7'h5 == reqIndex ? way0V_5 : _GEN_145; // @[DCache.scala 124:{33,33}]
  wire  _GEN_147 = 7'h6 == reqIndex ? way0V_6 : _GEN_146; // @[DCache.scala 124:{33,33}]
  wire  _GEN_148 = 7'h7 == reqIndex ? way0V_7 : _GEN_147; // @[DCache.scala 124:{33,33}]
  wire  _GEN_149 = 7'h8 == reqIndex ? way0V_8 : _GEN_148; // @[DCache.scala 124:{33,33}]
  wire  _GEN_150 = 7'h9 == reqIndex ? way0V_9 : _GEN_149; // @[DCache.scala 124:{33,33}]
  wire  _GEN_151 = 7'ha == reqIndex ? way0V_10 : _GEN_150; // @[DCache.scala 124:{33,33}]
  wire  _GEN_152 = 7'hb == reqIndex ? way0V_11 : _GEN_151; // @[DCache.scala 124:{33,33}]
  wire  _GEN_153 = 7'hc == reqIndex ? way0V_12 : _GEN_152; // @[DCache.scala 124:{33,33}]
  wire  _GEN_154 = 7'hd == reqIndex ? way0V_13 : _GEN_153; // @[DCache.scala 124:{33,33}]
  wire  _GEN_155 = 7'he == reqIndex ? way0V_14 : _GEN_154; // @[DCache.scala 124:{33,33}]
  wire  _GEN_156 = 7'hf == reqIndex ? way0V_15 : _GEN_155; // @[DCache.scala 124:{33,33}]
  wire  _GEN_157 = 7'h10 == reqIndex ? way0V_16 : _GEN_156; // @[DCache.scala 124:{33,33}]
  wire  _GEN_158 = 7'h11 == reqIndex ? way0V_17 : _GEN_157; // @[DCache.scala 124:{33,33}]
  wire  _GEN_159 = 7'h12 == reqIndex ? way0V_18 : _GEN_158; // @[DCache.scala 124:{33,33}]
  wire  _GEN_160 = 7'h13 == reqIndex ? way0V_19 : _GEN_159; // @[DCache.scala 124:{33,33}]
  wire  _GEN_161 = 7'h14 == reqIndex ? way0V_20 : _GEN_160; // @[DCache.scala 124:{33,33}]
  wire  _GEN_162 = 7'h15 == reqIndex ? way0V_21 : _GEN_161; // @[DCache.scala 124:{33,33}]
  wire  _GEN_163 = 7'h16 == reqIndex ? way0V_22 : _GEN_162; // @[DCache.scala 124:{33,33}]
  wire  _GEN_164 = 7'h17 == reqIndex ? way0V_23 : _GEN_163; // @[DCache.scala 124:{33,33}]
  wire  _GEN_165 = 7'h18 == reqIndex ? way0V_24 : _GEN_164; // @[DCache.scala 124:{33,33}]
  wire  _GEN_166 = 7'h19 == reqIndex ? way0V_25 : _GEN_165; // @[DCache.scala 124:{33,33}]
  wire  _GEN_167 = 7'h1a == reqIndex ? way0V_26 : _GEN_166; // @[DCache.scala 124:{33,33}]
  wire  _GEN_168 = 7'h1b == reqIndex ? way0V_27 : _GEN_167; // @[DCache.scala 124:{33,33}]
  wire  _GEN_169 = 7'h1c == reqIndex ? way0V_28 : _GEN_168; // @[DCache.scala 124:{33,33}]
  wire  _GEN_170 = 7'h1d == reqIndex ? way0V_29 : _GEN_169; // @[DCache.scala 124:{33,33}]
  wire  _GEN_171 = 7'h1e == reqIndex ? way0V_30 : _GEN_170; // @[DCache.scala 124:{33,33}]
  wire  _GEN_172 = 7'h1f == reqIndex ? way0V_31 : _GEN_171; // @[DCache.scala 124:{33,33}]
  wire  _GEN_173 = 7'h20 == reqIndex ? way0V_32 : _GEN_172; // @[DCache.scala 124:{33,33}]
  wire  _GEN_174 = 7'h21 == reqIndex ? way0V_33 : _GEN_173; // @[DCache.scala 124:{33,33}]
  wire  _GEN_175 = 7'h22 == reqIndex ? way0V_34 : _GEN_174; // @[DCache.scala 124:{33,33}]
  wire  _GEN_176 = 7'h23 == reqIndex ? way0V_35 : _GEN_175; // @[DCache.scala 124:{33,33}]
  wire  _GEN_177 = 7'h24 == reqIndex ? way0V_36 : _GEN_176; // @[DCache.scala 124:{33,33}]
  wire  _GEN_178 = 7'h25 == reqIndex ? way0V_37 : _GEN_177; // @[DCache.scala 124:{33,33}]
  wire  _GEN_179 = 7'h26 == reqIndex ? way0V_38 : _GEN_178; // @[DCache.scala 124:{33,33}]
  wire  _GEN_180 = 7'h27 == reqIndex ? way0V_39 : _GEN_179; // @[DCache.scala 124:{33,33}]
  wire  _GEN_181 = 7'h28 == reqIndex ? way0V_40 : _GEN_180; // @[DCache.scala 124:{33,33}]
  wire  _GEN_182 = 7'h29 == reqIndex ? way0V_41 : _GEN_181; // @[DCache.scala 124:{33,33}]
  wire  _GEN_183 = 7'h2a == reqIndex ? way0V_42 : _GEN_182; // @[DCache.scala 124:{33,33}]
  wire  _GEN_184 = 7'h2b == reqIndex ? way0V_43 : _GEN_183; // @[DCache.scala 124:{33,33}]
  wire  _GEN_185 = 7'h2c == reqIndex ? way0V_44 : _GEN_184; // @[DCache.scala 124:{33,33}]
  wire  _GEN_186 = 7'h2d == reqIndex ? way0V_45 : _GEN_185; // @[DCache.scala 124:{33,33}]
  wire  _GEN_187 = 7'h2e == reqIndex ? way0V_46 : _GEN_186; // @[DCache.scala 124:{33,33}]
  wire  _GEN_188 = 7'h2f == reqIndex ? way0V_47 : _GEN_187; // @[DCache.scala 124:{33,33}]
  wire  _GEN_189 = 7'h30 == reqIndex ? way0V_48 : _GEN_188; // @[DCache.scala 124:{33,33}]
  wire  _GEN_190 = 7'h31 == reqIndex ? way0V_49 : _GEN_189; // @[DCache.scala 124:{33,33}]
  wire  _GEN_191 = 7'h32 == reqIndex ? way0V_50 : _GEN_190; // @[DCache.scala 124:{33,33}]
  wire  _GEN_192 = 7'h33 == reqIndex ? way0V_51 : _GEN_191; // @[DCache.scala 124:{33,33}]
  wire  _GEN_193 = 7'h34 == reqIndex ? way0V_52 : _GEN_192; // @[DCache.scala 124:{33,33}]
  wire  _GEN_194 = 7'h35 == reqIndex ? way0V_53 : _GEN_193; // @[DCache.scala 124:{33,33}]
  wire  _GEN_195 = 7'h36 == reqIndex ? way0V_54 : _GEN_194; // @[DCache.scala 124:{33,33}]
  wire  _GEN_196 = 7'h37 == reqIndex ? way0V_55 : _GEN_195; // @[DCache.scala 124:{33,33}]
  wire  _GEN_197 = 7'h38 == reqIndex ? way0V_56 : _GEN_196; // @[DCache.scala 124:{33,33}]
  wire  _GEN_198 = 7'h39 == reqIndex ? way0V_57 : _GEN_197; // @[DCache.scala 124:{33,33}]
  wire  _GEN_199 = 7'h3a == reqIndex ? way0V_58 : _GEN_198; // @[DCache.scala 124:{33,33}]
  wire  _GEN_200 = 7'h3b == reqIndex ? way0V_59 : _GEN_199; // @[DCache.scala 124:{33,33}]
  wire  _GEN_201 = 7'h3c == reqIndex ? way0V_60 : _GEN_200; // @[DCache.scala 124:{33,33}]
  wire  _GEN_202 = 7'h3d == reqIndex ? way0V_61 : _GEN_201; // @[DCache.scala 124:{33,33}]
  wire  _GEN_203 = 7'h3e == reqIndex ? way0V_62 : _GEN_202; // @[DCache.scala 124:{33,33}]
  wire  _GEN_204 = 7'h3f == reqIndex ? way0V_63 : _GEN_203; // @[DCache.scala 124:{33,33}]
  wire  _GEN_205 = 7'h40 == reqIndex ? way0V_64 : _GEN_204; // @[DCache.scala 124:{33,33}]
  wire  _GEN_206 = 7'h41 == reqIndex ? way0V_65 : _GEN_205; // @[DCache.scala 124:{33,33}]
  wire  _GEN_207 = 7'h42 == reqIndex ? way0V_66 : _GEN_206; // @[DCache.scala 124:{33,33}]
  wire  _GEN_208 = 7'h43 == reqIndex ? way0V_67 : _GEN_207; // @[DCache.scala 124:{33,33}]
  wire  _GEN_209 = 7'h44 == reqIndex ? way0V_68 : _GEN_208; // @[DCache.scala 124:{33,33}]
  wire  _GEN_210 = 7'h45 == reqIndex ? way0V_69 : _GEN_209; // @[DCache.scala 124:{33,33}]
  wire  _GEN_211 = 7'h46 == reqIndex ? way0V_70 : _GEN_210; // @[DCache.scala 124:{33,33}]
  wire  _GEN_212 = 7'h47 == reqIndex ? way0V_71 : _GEN_211; // @[DCache.scala 124:{33,33}]
  wire  _GEN_213 = 7'h48 == reqIndex ? way0V_72 : _GEN_212; // @[DCache.scala 124:{33,33}]
  wire  _GEN_214 = 7'h49 == reqIndex ? way0V_73 : _GEN_213; // @[DCache.scala 124:{33,33}]
  wire  _GEN_215 = 7'h4a == reqIndex ? way0V_74 : _GEN_214; // @[DCache.scala 124:{33,33}]
  wire  _GEN_216 = 7'h4b == reqIndex ? way0V_75 : _GEN_215; // @[DCache.scala 124:{33,33}]
  wire  _GEN_217 = 7'h4c == reqIndex ? way0V_76 : _GEN_216; // @[DCache.scala 124:{33,33}]
  wire  _GEN_218 = 7'h4d == reqIndex ? way0V_77 : _GEN_217; // @[DCache.scala 124:{33,33}]
  wire  _GEN_219 = 7'h4e == reqIndex ? way0V_78 : _GEN_218; // @[DCache.scala 124:{33,33}]
  wire  _GEN_220 = 7'h4f == reqIndex ? way0V_79 : _GEN_219; // @[DCache.scala 124:{33,33}]
  wire  _GEN_221 = 7'h50 == reqIndex ? way0V_80 : _GEN_220; // @[DCache.scala 124:{33,33}]
  wire  _GEN_222 = 7'h51 == reqIndex ? way0V_81 : _GEN_221; // @[DCache.scala 124:{33,33}]
  wire  _GEN_223 = 7'h52 == reqIndex ? way0V_82 : _GEN_222; // @[DCache.scala 124:{33,33}]
  wire  _GEN_224 = 7'h53 == reqIndex ? way0V_83 : _GEN_223; // @[DCache.scala 124:{33,33}]
  wire  _GEN_225 = 7'h54 == reqIndex ? way0V_84 : _GEN_224; // @[DCache.scala 124:{33,33}]
  wire  _GEN_226 = 7'h55 == reqIndex ? way0V_85 : _GEN_225; // @[DCache.scala 124:{33,33}]
  wire  _GEN_227 = 7'h56 == reqIndex ? way0V_86 : _GEN_226; // @[DCache.scala 124:{33,33}]
  wire  _GEN_228 = 7'h57 == reqIndex ? way0V_87 : _GEN_227; // @[DCache.scala 124:{33,33}]
  wire  _GEN_229 = 7'h58 == reqIndex ? way0V_88 : _GEN_228; // @[DCache.scala 124:{33,33}]
  wire  _GEN_230 = 7'h59 == reqIndex ? way0V_89 : _GEN_229; // @[DCache.scala 124:{33,33}]
  wire  _GEN_231 = 7'h5a == reqIndex ? way0V_90 : _GEN_230; // @[DCache.scala 124:{33,33}]
  wire  _GEN_232 = 7'h5b == reqIndex ? way0V_91 : _GEN_231; // @[DCache.scala 124:{33,33}]
  wire  _GEN_233 = 7'h5c == reqIndex ? way0V_92 : _GEN_232; // @[DCache.scala 124:{33,33}]
  wire  _GEN_234 = 7'h5d == reqIndex ? way0V_93 : _GEN_233; // @[DCache.scala 124:{33,33}]
  wire  _GEN_235 = 7'h5e == reqIndex ? way0V_94 : _GEN_234; // @[DCache.scala 124:{33,33}]
  wire  _GEN_236 = 7'h5f == reqIndex ? way0V_95 : _GEN_235; // @[DCache.scala 124:{33,33}]
  wire  _GEN_237 = 7'h60 == reqIndex ? way0V_96 : _GEN_236; // @[DCache.scala 124:{33,33}]
  wire  _GEN_238 = 7'h61 == reqIndex ? way0V_97 : _GEN_237; // @[DCache.scala 124:{33,33}]
  wire  _GEN_239 = 7'h62 == reqIndex ? way0V_98 : _GEN_238; // @[DCache.scala 124:{33,33}]
  wire  _GEN_240 = 7'h63 == reqIndex ? way0V_99 : _GEN_239; // @[DCache.scala 124:{33,33}]
  wire  _GEN_241 = 7'h64 == reqIndex ? way0V_100 : _GEN_240; // @[DCache.scala 124:{33,33}]
  wire  _GEN_242 = 7'h65 == reqIndex ? way0V_101 : _GEN_241; // @[DCache.scala 124:{33,33}]
  wire  _GEN_243 = 7'h66 == reqIndex ? way0V_102 : _GEN_242; // @[DCache.scala 124:{33,33}]
  wire  _GEN_244 = 7'h67 == reqIndex ? way0V_103 : _GEN_243; // @[DCache.scala 124:{33,33}]
  wire  _GEN_245 = 7'h68 == reqIndex ? way0V_104 : _GEN_244; // @[DCache.scala 124:{33,33}]
  wire  _GEN_246 = 7'h69 == reqIndex ? way0V_105 : _GEN_245; // @[DCache.scala 124:{33,33}]
  wire  _GEN_247 = 7'h6a == reqIndex ? way0V_106 : _GEN_246; // @[DCache.scala 124:{33,33}]
  wire  _GEN_248 = 7'h6b == reqIndex ? way0V_107 : _GEN_247; // @[DCache.scala 124:{33,33}]
  wire  _GEN_249 = 7'h6c == reqIndex ? way0V_108 : _GEN_248; // @[DCache.scala 124:{33,33}]
  wire  _GEN_250 = 7'h6d == reqIndex ? way0V_109 : _GEN_249; // @[DCache.scala 124:{33,33}]
  wire  _GEN_251 = 7'h6e == reqIndex ? way0V_110 : _GEN_250; // @[DCache.scala 124:{33,33}]
  wire  _GEN_252 = 7'h6f == reqIndex ? way0V_111 : _GEN_251; // @[DCache.scala 124:{33,33}]
  wire  _GEN_253 = 7'h70 == reqIndex ? way0V_112 : _GEN_252; // @[DCache.scala 124:{33,33}]
  wire  _GEN_254 = 7'h71 == reqIndex ? way0V_113 : _GEN_253; // @[DCache.scala 124:{33,33}]
  wire  _GEN_255 = 7'h72 == reqIndex ? way0V_114 : _GEN_254; // @[DCache.scala 124:{33,33}]
  wire  _GEN_256 = 7'h73 == reqIndex ? way0V_115 : _GEN_255; // @[DCache.scala 124:{33,33}]
  wire  _GEN_257 = 7'h74 == reqIndex ? way0V_116 : _GEN_256; // @[DCache.scala 124:{33,33}]
  wire  _GEN_258 = 7'h75 == reqIndex ? way0V_117 : _GEN_257; // @[DCache.scala 124:{33,33}]
  wire  _GEN_259 = 7'h76 == reqIndex ? way0V_118 : _GEN_258; // @[DCache.scala 124:{33,33}]
  wire  _GEN_260 = 7'h77 == reqIndex ? way0V_119 : _GEN_259; // @[DCache.scala 124:{33,33}]
  wire  _GEN_261 = 7'h78 == reqIndex ? way0V_120 : _GEN_260; // @[DCache.scala 124:{33,33}]
  wire  _GEN_262 = 7'h79 == reqIndex ? way0V_121 : _GEN_261; // @[DCache.scala 124:{33,33}]
  wire  _GEN_263 = 7'h7a == reqIndex ? way0V_122 : _GEN_262; // @[DCache.scala 124:{33,33}]
  wire  _GEN_264 = 7'h7b == reqIndex ? way0V_123 : _GEN_263; // @[DCache.scala 124:{33,33}]
  wire  _GEN_265 = 7'h7c == reqIndex ? way0V_124 : _GEN_264; // @[DCache.scala 124:{33,33}]
  wire  _GEN_266 = 7'h7d == reqIndex ? way0V_125 : _GEN_265; // @[DCache.scala 124:{33,33}]
  wire  _GEN_267 = 7'h7e == reqIndex ? way0V_126 : _GEN_266; // @[DCache.scala 124:{33,33}]
  wire  _GEN_268 = 7'h7f == reqIndex ? way0V_127 : _GEN_267; // @[DCache.scala 124:{33,33}]
  wire [20:0] _GEN_14 = 7'h1 == reqIndex ? way0Tag_1 : way0Tag_0; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_15 = 7'h2 == reqIndex ? way0Tag_2 : _GEN_14; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_16 = 7'h3 == reqIndex ? way0Tag_3 : _GEN_15; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_17 = 7'h4 == reqIndex ? way0Tag_4 : _GEN_16; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_18 = 7'h5 == reqIndex ? way0Tag_5 : _GEN_17; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_19 = 7'h6 == reqIndex ? way0Tag_6 : _GEN_18; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_20 = 7'h7 == reqIndex ? way0Tag_7 : _GEN_19; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_21 = 7'h8 == reqIndex ? way0Tag_8 : _GEN_20; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_22 = 7'h9 == reqIndex ? way0Tag_9 : _GEN_21; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_23 = 7'ha == reqIndex ? way0Tag_10 : _GEN_22; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_24 = 7'hb == reqIndex ? way0Tag_11 : _GEN_23; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_25 = 7'hc == reqIndex ? way0Tag_12 : _GEN_24; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_26 = 7'hd == reqIndex ? way0Tag_13 : _GEN_25; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_27 = 7'he == reqIndex ? way0Tag_14 : _GEN_26; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_28 = 7'hf == reqIndex ? way0Tag_15 : _GEN_27; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_29 = 7'h10 == reqIndex ? way0Tag_16 : _GEN_28; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_30 = 7'h11 == reqIndex ? way0Tag_17 : _GEN_29; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_31 = 7'h12 == reqIndex ? way0Tag_18 : _GEN_30; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_32 = 7'h13 == reqIndex ? way0Tag_19 : _GEN_31; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_33 = 7'h14 == reqIndex ? way0Tag_20 : _GEN_32; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_34 = 7'h15 == reqIndex ? way0Tag_21 : _GEN_33; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_35 = 7'h16 == reqIndex ? way0Tag_22 : _GEN_34; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_36 = 7'h17 == reqIndex ? way0Tag_23 : _GEN_35; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_37 = 7'h18 == reqIndex ? way0Tag_24 : _GEN_36; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_38 = 7'h19 == reqIndex ? way0Tag_25 : _GEN_37; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_39 = 7'h1a == reqIndex ? way0Tag_26 : _GEN_38; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_40 = 7'h1b == reqIndex ? way0Tag_27 : _GEN_39; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_41 = 7'h1c == reqIndex ? way0Tag_28 : _GEN_40; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_42 = 7'h1d == reqIndex ? way0Tag_29 : _GEN_41; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_43 = 7'h1e == reqIndex ? way0Tag_30 : _GEN_42; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_44 = 7'h1f == reqIndex ? way0Tag_31 : _GEN_43; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_45 = 7'h20 == reqIndex ? way0Tag_32 : _GEN_44; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_46 = 7'h21 == reqIndex ? way0Tag_33 : _GEN_45; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_47 = 7'h22 == reqIndex ? way0Tag_34 : _GEN_46; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_48 = 7'h23 == reqIndex ? way0Tag_35 : _GEN_47; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_49 = 7'h24 == reqIndex ? way0Tag_36 : _GEN_48; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_50 = 7'h25 == reqIndex ? way0Tag_37 : _GEN_49; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_51 = 7'h26 == reqIndex ? way0Tag_38 : _GEN_50; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_52 = 7'h27 == reqIndex ? way0Tag_39 : _GEN_51; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_53 = 7'h28 == reqIndex ? way0Tag_40 : _GEN_52; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_54 = 7'h29 == reqIndex ? way0Tag_41 : _GEN_53; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_55 = 7'h2a == reqIndex ? way0Tag_42 : _GEN_54; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_56 = 7'h2b == reqIndex ? way0Tag_43 : _GEN_55; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_57 = 7'h2c == reqIndex ? way0Tag_44 : _GEN_56; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_58 = 7'h2d == reqIndex ? way0Tag_45 : _GEN_57; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_59 = 7'h2e == reqIndex ? way0Tag_46 : _GEN_58; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_60 = 7'h2f == reqIndex ? way0Tag_47 : _GEN_59; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_61 = 7'h30 == reqIndex ? way0Tag_48 : _GEN_60; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_62 = 7'h31 == reqIndex ? way0Tag_49 : _GEN_61; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_63 = 7'h32 == reqIndex ? way0Tag_50 : _GEN_62; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_64 = 7'h33 == reqIndex ? way0Tag_51 : _GEN_63; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_65 = 7'h34 == reqIndex ? way0Tag_52 : _GEN_64; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_66 = 7'h35 == reqIndex ? way0Tag_53 : _GEN_65; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_67 = 7'h36 == reqIndex ? way0Tag_54 : _GEN_66; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_68 = 7'h37 == reqIndex ? way0Tag_55 : _GEN_67; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_69 = 7'h38 == reqIndex ? way0Tag_56 : _GEN_68; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_70 = 7'h39 == reqIndex ? way0Tag_57 : _GEN_69; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_71 = 7'h3a == reqIndex ? way0Tag_58 : _GEN_70; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_72 = 7'h3b == reqIndex ? way0Tag_59 : _GEN_71; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_73 = 7'h3c == reqIndex ? way0Tag_60 : _GEN_72; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_74 = 7'h3d == reqIndex ? way0Tag_61 : _GEN_73; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_75 = 7'h3e == reqIndex ? way0Tag_62 : _GEN_74; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_76 = 7'h3f == reqIndex ? way0Tag_63 : _GEN_75; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_77 = 7'h40 == reqIndex ? way0Tag_64 : _GEN_76; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_78 = 7'h41 == reqIndex ? way0Tag_65 : _GEN_77; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_79 = 7'h42 == reqIndex ? way0Tag_66 : _GEN_78; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_80 = 7'h43 == reqIndex ? way0Tag_67 : _GEN_79; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_81 = 7'h44 == reqIndex ? way0Tag_68 : _GEN_80; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_82 = 7'h45 == reqIndex ? way0Tag_69 : _GEN_81; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_83 = 7'h46 == reqIndex ? way0Tag_70 : _GEN_82; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_84 = 7'h47 == reqIndex ? way0Tag_71 : _GEN_83; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_85 = 7'h48 == reqIndex ? way0Tag_72 : _GEN_84; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_86 = 7'h49 == reqIndex ? way0Tag_73 : _GEN_85; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_87 = 7'h4a == reqIndex ? way0Tag_74 : _GEN_86; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_88 = 7'h4b == reqIndex ? way0Tag_75 : _GEN_87; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_89 = 7'h4c == reqIndex ? way0Tag_76 : _GEN_88; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_90 = 7'h4d == reqIndex ? way0Tag_77 : _GEN_89; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_91 = 7'h4e == reqIndex ? way0Tag_78 : _GEN_90; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_92 = 7'h4f == reqIndex ? way0Tag_79 : _GEN_91; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_93 = 7'h50 == reqIndex ? way0Tag_80 : _GEN_92; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_94 = 7'h51 == reqIndex ? way0Tag_81 : _GEN_93; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_95 = 7'h52 == reqIndex ? way0Tag_82 : _GEN_94; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_96 = 7'h53 == reqIndex ? way0Tag_83 : _GEN_95; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_97 = 7'h54 == reqIndex ? way0Tag_84 : _GEN_96; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_98 = 7'h55 == reqIndex ? way0Tag_85 : _GEN_97; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_99 = 7'h56 == reqIndex ? way0Tag_86 : _GEN_98; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_100 = 7'h57 == reqIndex ? way0Tag_87 : _GEN_99; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_101 = 7'h58 == reqIndex ? way0Tag_88 : _GEN_100; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_102 = 7'h59 == reqIndex ? way0Tag_89 : _GEN_101; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_103 = 7'h5a == reqIndex ? way0Tag_90 : _GEN_102; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_104 = 7'h5b == reqIndex ? way0Tag_91 : _GEN_103; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_105 = 7'h5c == reqIndex ? way0Tag_92 : _GEN_104; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_106 = 7'h5d == reqIndex ? way0Tag_93 : _GEN_105; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_107 = 7'h5e == reqIndex ? way0Tag_94 : _GEN_106; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_108 = 7'h5f == reqIndex ? way0Tag_95 : _GEN_107; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_109 = 7'h60 == reqIndex ? way0Tag_96 : _GEN_108; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_110 = 7'h61 == reqIndex ? way0Tag_97 : _GEN_109; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_111 = 7'h62 == reqIndex ? way0Tag_98 : _GEN_110; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_112 = 7'h63 == reqIndex ? way0Tag_99 : _GEN_111; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_113 = 7'h64 == reqIndex ? way0Tag_100 : _GEN_112; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_114 = 7'h65 == reqIndex ? way0Tag_101 : _GEN_113; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_115 = 7'h66 == reqIndex ? way0Tag_102 : _GEN_114; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_116 = 7'h67 == reqIndex ? way0Tag_103 : _GEN_115; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_117 = 7'h68 == reqIndex ? way0Tag_104 : _GEN_116; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_118 = 7'h69 == reqIndex ? way0Tag_105 : _GEN_117; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_119 = 7'h6a == reqIndex ? way0Tag_106 : _GEN_118; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_120 = 7'h6b == reqIndex ? way0Tag_107 : _GEN_119; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_121 = 7'h6c == reqIndex ? way0Tag_108 : _GEN_120; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_122 = 7'h6d == reqIndex ? way0Tag_109 : _GEN_121; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_123 = 7'h6e == reqIndex ? way0Tag_110 : _GEN_122; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_124 = 7'h6f == reqIndex ? way0Tag_111 : _GEN_123; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_125 = 7'h70 == reqIndex ? way0Tag_112 : _GEN_124; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_126 = 7'h71 == reqIndex ? way0Tag_113 : _GEN_125; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_127 = 7'h72 == reqIndex ? way0Tag_114 : _GEN_126; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_128 = 7'h73 == reqIndex ? way0Tag_115 : _GEN_127; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_129 = 7'h74 == reqIndex ? way0Tag_116 : _GEN_128; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_130 = 7'h75 == reqIndex ? way0Tag_117 : _GEN_129; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_131 = 7'h76 == reqIndex ? way0Tag_118 : _GEN_130; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_132 = 7'h77 == reqIndex ? way0Tag_119 : _GEN_131; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_133 = 7'h78 == reqIndex ? way0Tag_120 : _GEN_132; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_134 = 7'h79 == reqIndex ? way0Tag_121 : _GEN_133; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_135 = 7'h7a == reqIndex ? way0Tag_122 : _GEN_134; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_136 = 7'h7b == reqIndex ? way0Tag_123 : _GEN_135; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_137 = 7'h7c == reqIndex ? way0Tag_124 : _GEN_136; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_138 = 7'h7d == reqIndex ? way0Tag_125 : _GEN_137; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_139 = 7'h7e == reqIndex ? way0Tag_126 : _GEN_138; // @[DCache.scala 124:{55,55}]
  wire [20:0] _GEN_140 = 7'h7f == reqIndex ? way0Tag_127 : _GEN_139; // @[DCache.scala 124:{55,55}]
  wire  way0Hit = _GEN_268 & _GEN_140 == reqTag; // @[DCache.scala 124:33]
  wire  _GEN_398 = 7'h1 == reqIndex ? way1V_1 : way1V_0; // @[DCache.scala 125:{33,33}]
  wire  _GEN_399 = 7'h2 == reqIndex ? way1V_2 : _GEN_398; // @[DCache.scala 125:{33,33}]
  wire  _GEN_400 = 7'h3 == reqIndex ? way1V_3 : _GEN_399; // @[DCache.scala 125:{33,33}]
  wire  _GEN_401 = 7'h4 == reqIndex ? way1V_4 : _GEN_400; // @[DCache.scala 125:{33,33}]
  wire  _GEN_402 = 7'h5 == reqIndex ? way1V_5 : _GEN_401; // @[DCache.scala 125:{33,33}]
  wire  _GEN_403 = 7'h6 == reqIndex ? way1V_6 : _GEN_402; // @[DCache.scala 125:{33,33}]
  wire  _GEN_404 = 7'h7 == reqIndex ? way1V_7 : _GEN_403; // @[DCache.scala 125:{33,33}]
  wire  _GEN_405 = 7'h8 == reqIndex ? way1V_8 : _GEN_404; // @[DCache.scala 125:{33,33}]
  wire  _GEN_406 = 7'h9 == reqIndex ? way1V_9 : _GEN_405; // @[DCache.scala 125:{33,33}]
  wire  _GEN_407 = 7'ha == reqIndex ? way1V_10 : _GEN_406; // @[DCache.scala 125:{33,33}]
  wire  _GEN_408 = 7'hb == reqIndex ? way1V_11 : _GEN_407; // @[DCache.scala 125:{33,33}]
  wire  _GEN_409 = 7'hc == reqIndex ? way1V_12 : _GEN_408; // @[DCache.scala 125:{33,33}]
  wire  _GEN_410 = 7'hd == reqIndex ? way1V_13 : _GEN_409; // @[DCache.scala 125:{33,33}]
  wire  _GEN_411 = 7'he == reqIndex ? way1V_14 : _GEN_410; // @[DCache.scala 125:{33,33}]
  wire  _GEN_412 = 7'hf == reqIndex ? way1V_15 : _GEN_411; // @[DCache.scala 125:{33,33}]
  wire  _GEN_413 = 7'h10 == reqIndex ? way1V_16 : _GEN_412; // @[DCache.scala 125:{33,33}]
  wire  _GEN_414 = 7'h11 == reqIndex ? way1V_17 : _GEN_413; // @[DCache.scala 125:{33,33}]
  wire  _GEN_415 = 7'h12 == reqIndex ? way1V_18 : _GEN_414; // @[DCache.scala 125:{33,33}]
  wire  _GEN_416 = 7'h13 == reqIndex ? way1V_19 : _GEN_415; // @[DCache.scala 125:{33,33}]
  wire  _GEN_417 = 7'h14 == reqIndex ? way1V_20 : _GEN_416; // @[DCache.scala 125:{33,33}]
  wire  _GEN_418 = 7'h15 == reqIndex ? way1V_21 : _GEN_417; // @[DCache.scala 125:{33,33}]
  wire  _GEN_419 = 7'h16 == reqIndex ? way1V_22 : _GEN_418; // @[DCache.scala 125:{33,33}]
  wire  _GEN_420 = 7'h17 == reqIndex ? way1V_23 : _GEN_419; // @[DCache.scala 125:{33,33}]
  wire  _GEN_421 = 7'h18 == reqIndex ? way1V_24 : _GEN_420; // @[DCache.scala 125:{33,33}]
  wire  _GEN_422 = 7'h19 == reqIndex ? way1V_25 : _GEN_421; // @[DCache.scala 125:{33,33}]
  wire  _GEN_423 = 7'h1a == reqIndex ? way1V_26 : _GEN_422; // @[DCache.scala 125:{33,33}]
  wire  _GEN_424 = 7'h1b == reqIndex ? way1V_27 : _GEN_423; // @[DCache.scala 125:{33,33}]
  wire  _GEN_425 = 7'h1c == reqIndex ? way1V_28 : _GEN_424; // @[DCache.scala 125:{33,33}]
  wire  _GEN_426 = 7'h1d == reqIndex ? way1V_29 : _GEN_425; // @[DCache.scala 125:{33,33}]
  wire  _GEN_427 = 7'h1e == reqIndex ? way1V_30 : _GEN_426; // @[DCache.scala 125:{33,33}]
  wire  _GEN_428 = 7'h1f == reqIndex ? way1V_31 : _GEN_427; // @[DCache.scala 125:{33,33}]
  wire  _GEN_429 = 7'h20 == reqIndex ? way1V_32 : _GEN_428; // @[DCache.scala 125:{33,33}]
  wire  _GEN_430 = 7'h21 == reqIndex ? way1V_33 : _GEN_429; // @[DCache.scala 125:{33,33}]
  wire  _GEN_431 = 7'h22 == reqIndex ? way1V_34 : _GEN_430; // @[DCache.scala 125:{33,33}]
  wire  _GEN_432 = 7'h23 == reqIndex ? way1V_35 : _GEN_431; // @[DCache.scala 125:{33,33}]
  wire  _GEN_433 = 7'h24 == reqIndex ? way1V_36 : _GEN_432; // @[DCache.scala 125:{33,33}]
  wire  _GEN_434 = 7'h25 == reqIndex ? way1V_37 : _GEN_433; // @[DCache.scala 125:{33,33}]
  wire  _GEN_435 = 7'h26 == reqIndex ? way1V_38 : _GEN_434; // @[DCache.scala 125:{33,33}]
  wire  _GEN_436 = 7'h27 == reqIndex ? way1V_39 : _GEN_435; // @[DCache.scala 125:{33,33}]
  wire  _GEN_437 = 7'h28 == reqIndex ? way1V_40 : _GEN_436; // @[DCache.scala 125:{33,33}]
  wire  _GEN_438 = 7'h29 == reqIndex ? way1V_41 : _GEN_437; // @[DCache.scala 125:{33,33}]
  wire  _GEN_439 = 7'h2a == reqIndex ? way1V_42 : _GEN_438; // @[DCache.scala 125:{33,33}]
  wire  _GEN_440 = 7'h2b == reqIndex ? way1V_43 : _GEN_439; // @[DCache.scala 125:{33,33}]
  wire  _GEN_441 = 7'h2c == reqIndex ? way1V_44 : _GEN_440; // @[DCache.scala 125:{33,33}]
  wire  _GEN_442 = 7'h2d == reqIndex ? way1V_45 : _GEN_441; // @[DCache.scala 125:{33,33}]
  wire  _GEN_443 = 7'h2e == reqIndex ? way1V_46 : _GEN_442; // @[DCache.scala 125:{33,33}]
  wire  _GEN_444 = 7'h2f == reqIndex ? way1V_47 : _GEN_443; // @[DCache.scala 125:{33,33}]
  wire  _GEN_445 = 7'h30 == reqIndex ? way1V_48 : _GEN_444; // @[DCache.scala 125:{33,33}]
  wire  _GEN_446 = 7'h31 == reqIndex ? way1V_49 : _GEN_445; // @[DCache.scala 125:{33,33}]
  wire  _GEN_447 = 7'h32 == reqIndex ? way1V_50 : _GEN_446; // @[DCache.scala 125:{33,33}]
  wire  _GEN_448 = 7'h33 == reqIndex ? way1V_51 : _GEN_447; // @[DCache.scala 125:{33,33}]
  wire  _GEN_449 = 7'h34 == reqIndex ? way1V_52 : _GEN_448; // @[DCache.scala 125:{33,33}]
  wire  _GEN_450 = 7'h35 == reqIndex ? way1V_53 : _GEN_449; // @[DCache.scala 125:{33,33}]
  wire  _GEN_451 = 7'h36 == reqIndex ? way1V_54 : _GEN_450; // @[DCache.scala 125:{33,33}]
  wire  _GEN_452 = 7'h37 == reqIndex ? way1V_55 : _GEN_451; // @[DCache.scala 125:{33,33}]
  wire  _GEN_453 = 7'h38 == reqIndex ? way1V_56 : _GEN_452; // @[DCache.scala 125:{33,33}]
  wire  _GEN_454 = 7'h39 == reqIndex ? way1V_57 : _GEN_453; // @[DCache.scala 125:{33,33}]
  wire  _GEN_455 = 7'h3a == reqIndex ? way1V_58 : _GEN_454; // @[DCache.scala 125:{33,33}]
  wire  _GEN_456 = 7'h3b == reqIndex ? way1V_59 : _GEN_455; // @[DCache.scala 125:{33,33}]
  wire  _GEN_457 = 7'h3c == reqIndex ? way1V_60 : _GEN_456; // @[DCache.scala 125:{33,33}]
  wire  _GEN_458 = 7'h3d == reqIndex ? way1V_61 : _GEN_457; // @[DCache.scala 125:{33,33}]
  wire  _GEN_459 = 7'h3e == reqIndex ? way1V_62 : _GEN_458; // @[DCache.scala 125:{33,33}]
  wire  _GEN_460 = 7'h3f == reqIndex ? way1V_63 : _GEN_459; // @[DCache.scala 125:{33,33}]
  wire  _GEN_461 = 7'h40 == reqIndex ? way1V_64 : _GEN_460; // @[DCache.scala 125:{33,33}]
  wire  _GEN_462 = 7'h41 == reqIndex ? way1V_65 : _GEN_461; // @[DCache.scala 125:{33,33}]
  wire  _GEN_463 = 7'h42 == reqIndex ? way1V_66 : _GEN_462; // @[DCache.scala 125:{33,33}]
  wire  _GEN_464 = 7'h43 == reqIndex ? way1V_67 : _GEN_463; // @[DCache.scala 125:{33,33}]
  wire  _GEN_465 = 7'h44 == reqIndex ? way1V_68 : _GEN_464; // @[DCache.scala 125:{33,33}]
  wire  _GEN_466 = 7'h45 == reqIndex ? way1V_69 : _GEN_465; // @[DCache.scala 125:{33,33}]
  wire  _GEN_467 = 7'h46 == reqIndex ? way1V_70 : _GEN_466; // @[DCache.scala 125:{33,33}]
  wire  _GEN_468 = 7'h47 == reqIndex ? way1V_71 : _GEN_467; // @[DCache.scala 125:{33,33}]
  wire  _GEN_469 = 7'h48 == reqIndex ? way1V_72 : _GEN_468; // @[DCache.scala 125:{33,33}]
  wire  _GEN_470 = 7'h49 == reqIndex ? way1V_73 : _GEN_469; // @[DCache.scala 125:{33,33}]
  wire  _GEN_471 = 7'h4a == reqIndex ? way1V_74 : _GEN_470; // @[DCache.scala 125:{33,33}]
  wire  _GEN_472 = 7'h4b == reqIndex ? way1V_75 : _GEN_471; // @[DCache.scala 125:{33,33}]
  wire  _GEN_473 = 7'h4c == reqIndex ? way1V_76 : _GEN_472; // @[DCache.scala 125:{33,33}]
  wire  _GEN_474 = 7'h4d == reqIndex ? way1V_77 : _GEN_473; // @[DCache.scala 125:{33,33}]
  wire  _GEN_475 = 7'h4e == reqIndex ? way1V_78 : _GEN_474; // @[DCache.scala 125:{33,33}]
  wire  _GEN_476 = 7'h4f == reqIndex ? way1V_79 : _GEN_475; // @[DCache.scala 125:{33,33}]
  wire  _GEN_477 = 7'h50 == reqIndex ? way1V_80 : _GEN_476; // @[DCache.scala 125:{33,33}]
  wire  _GEN_478 = 7'h51 == reqIndex ? way1V_81 : _GEN_477; // @[DCache.scala 125:{33,33}]
  wire  _GEN_479 = 7'h52 == reqIndex ? way1V_82 : _GEN_478; // @[DCache.scala 125:{33,33}]
  wire  _GEN_480 = 7'h53 == reqIndex ? way1V_83 : _GEN_479; // @[DCache.scala 125:{33,33}]
  wire  _GEN_481 = 7'h54 == reqIndex ? way1V_84 : _GEN_480; // @[DCache.scala 125:{33,33}]
  wire  _GEN_482 = 7'h55 == reqIndex ? way1V_85 : _GEN_481; // @[DCache.scala 125:{33,33}]
  wire  _GEN_483 = 7'h56 == reqIndex ? way1V_86 : _GEN_482; // @[DCache.scala 125:{33,33}]
  wire  _GEN_484 = 7'h57 == reqIndex ? way1V_87 : _GEN_483; // @[DCache.scala 125:{33,33}]
  wire  _GEN_485 = 7'h58 == reqIndex ? way1V_88 : _GEN_484; // @[DCache.scala 125:{33,33}]
  wire  _GEN_486 = 7'h59 == reqIndex ? way1V_89 : _GEN_485; // @[DCache.scala 125:{33,33}]
  wire  _GEN_487 = 7'h5a == reqIndex ? way1V_90 : _GEN_486; // @[DCache.scala 125:{33,33}]
  wire  _GEN_488 = 7'h5b == reqIndex ? way1V_91 : _GEN_487; // @[DCache.scala 125:{33,33}]
  wire  _GEN_489 = 7'h5c == reqIndex ? way1V_92 : _GEN_488; // @[DCache.scala 125:{33,33}]
  wire  _GEN_490 = 7'h5d == reqIndex ? way1V_93 : _GEN_489; // @[DCache.scala 125:{33,33}]
  wire  _GEN_491 = 7'h5e == reqIndex ? way1V_94 : _GEN_490; // @[DCache.scala 125:{33,33}]
  wire  _GEN_492 = 7'h5f == reqIndex ? way1V_95 : _GEN_491; // @[DCache.scala 125:{33,33}]
  wire  _GEN_493 = 7'h60 == reqIndex ? way1V_96 : _GEN_492; // @[DCache.scala 125:{33,33}]
  wire  _GEN_494 = 7'h61 == reqIndex ? way1V_97 : _GEN_493; // @[DCache.scala 125:{33,33}]
  wire  _GEN_495 = 7'h62 == reqIndex ? way1V_98 : _GEN_494; // @[DCache.scala 125:{33,33}]
  wire  _GEN_496 = 7'h63 == reqIndex ? way1V_99 : _GEN_495; // @[DCache.scala 125:{33,33}]
  wire  _GEN_497 = 7'h64 == reqIndex ? way1V_100 : _GEN_496; // @[DCache.scala 125:{33,33}]
  wire  _GEN_498 = 7'h65 == reqIndex ? way1V_101 : _GEN_497; // @[DCache.scala 125:{33,33}]
  wire  _GEN_499 = 7'h66 == reqIndex ? way1V_102 : _GEN_498; // @[DCache.scala 125:{33,33}]
  wire  _GEN_500 = 7'h67 == reqIndex ? way1V_103 : _GEN_499; // @[DCache.scala 125:{33,33}]
  wire  _GEN_501 = 7'h68 == reqIndex ? way1V_104 : _GEN_500; // @[DCache.scala 125:{33,33}]
  wire  _GEN_502 = 7'h69 == reqIndex ? way1V_105 : _GEN_501; // @[DCache.scala 125:{33,33}]
  wire  _GEN_503 = 7'h6a == reqIndex ? way1V_106 : _GEN_502; // @[DCache.scala 125:{33,33}]
  wire  _GEN_504 = 7'h6b == reqIndex ? way1V_107 : _GEN_503; // @[DCache.scala 125:{33,33}]
  wire  _GEN_505 = 7'h6c == reqIndex ? way1V_108 : _GEN_504; // @[DCache.scala 125:{33,33}]
  wire  _GEN_506 = 7'h6d == reqIndex ? way1V_109 : _GEN_505; // @[DCache.scala 125:{33,33}]
  wire  _GEN_507 = 7'h6e == reqIndex ? way1V_110 : _GEN_506; // @[DCache.scala 125:{33,33}]
  wire  _GEN_508 = 7'h6f == reqIndex ? way1V_111 : _GEN_507; // @[DCache.scala 125:{33,33}]
  wire  _GEN_509 = 7'h70 == reqIndex ? way1V_112 : _GEN_508; // @[DCache.scala 125:{33,33}]
  wire  _GEN_510 = 7'h71 == reqIndex ? way1V_113 : _GEN_509; // @[DCache.scala 125:{33,33}]
  wire  _GEN_511 = 7'h72 == reqIndex ? way1V_114 : _GEN_510; // @[DCache.scala 125:{33,33}]
  wire  _GEN_512 = 7'h73 == reqIndex ? way1V_115 : _GEN_511; // @[DCache.scala 125:{33,33}]
  wire  _GEN_513 = 7'h74 == reqIndex ? way1V_116 : _GEN_512; // @[DCache.scala 125:{33,33}]
  wire  _GEN_514 = 7'h75 == reqIndex ? way1V_117 : _GEN_513; // @[DCache.scala 125:{33,33}]
  wire  _GEN_515 = 7'h76 == reqIndex ? way1V_118 : _GEN_514; // @[DCache.scala 125:{33,33}]
  wire  _GEN_516 = 7'h77 == reqIndex ? way1V_119 : _GEN_515; // @[DCache.scala 125:{33,33}]
  wire  _GEN_517 = 7'h78 == reqIndex ? way1V_120 : _GEN_516; // @[DCache.scala 125:{33,33}]
  wire  _GEN_518 = 7'h79 == reqIndex ? way1V_121 : _GEN_517; // @[DCache.scala 125:{33,33}]
  wire  _GEN_519 = 7'h7a == reqIndex ? way1V_122 : _GEN_518; // @[DCache.scala 125:{33,33}]
  wire  _GEN_520 = 7'h7b == reqIndex ? way1V_123 : _GEN_519; // @[DCache.scala 125:{33,33}]
  wire  _GEN_521 = 7'h7c == reqIndex ? way1V_124 : _GEN_520; // @[DCache.scala 125:{33,33}]
  wire  _GEN_522 = 7'h7d == reqIndex ? way1V_125 : _GEN_521; // @[DCache.scala 125:{33,33}]
  wire  _GEN_523 = 7'h7e == reqIndex ? way1V_126 : _GEN_522; // @[DCache.scala 125:{33,33}]
  wire  _GEN_524 = 7'h7f == reqIndex ? way1V_127 : _GEN_523; // @[DCache.scala 125:{33,33}]
  wire [20:0] _GEN_270 = 7'h1 == reqIndex ? way1Tag_1 : way1Tag_0; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_271 = 7'h2 == reqIndex ? way1Tag_2 : _GEN_270; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_272 = 7'h3 == reqIndex ? way1Tag_3 : _GEN_271; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_273 = 7'h4 == reqIndex ? way1Tag_4 : _GEN_272; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_274 = 7'h5 == reqIndex ? way1Tag_5 : _GEN_273; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_275 = 7'h6 == reqIndex ? way1Tag_6 : _GEN_274; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_276 = 7'h7 == reqIndex ? way1Tag_7 : _GEN_275; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_277 = 7'h8 == reqIndex ? way1Tag_8 : _GEN_276; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_278 = 7'h9 == reqIndex ? way1Tag_9 : _GEN_277; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_279 = 7'ha == reqIndex ? way1Tag_10 : _GEN_278; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_280 = 7'hb == reqIndex ? way1Tag_11 : _GEN_279; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_281 = 7'hc == reqIndex ? way1Tag_12 : _GEN_280; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_282 = 7'hd == reqIndex ? way1Tag_13 : _GEN_281; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_283 = 7'he == reqIndex ? way1Tag_14 : _GEN_282; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_284 = 7'hf == reqIndex ? way1Tag_15 : _GEN_283; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_285 = 7'h10 == reqIndex ? way1Tag_16 : _GEN_284; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_286 = 7'h11 == reqIndex ? way1Tag_17 : _GEN_285; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_287 = 7'h12 == reqIndex ? way1Tag_18 : _GEN_286; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_288 = 7'h13 == reqIndex ? way1Tag_19 : _GEN_287; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_289 = 7'h14 == reqIndex ? way1Tag_20 : _GEN_288; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_290 = 7'h15 == reqIndex ? way1Tag_21 : _GEN_289; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_291 = 7'h16 == reqIndex ? way1Tag_22 : _GEN_290; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_292 = 7'h17 == reqIndex ? way1Tag_23 : _GEN_291; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_293 = 7'h18 == reqIndex ? way1Tag_24 : _GEN_292; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_294 = 7'h19 == reqIndex ? way1Tag_25 : _GEN_293; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_295 = 7'h1a == reqIndex ? way1Tag_26 : _GEN_294; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_296 = 7'h1b == reqIndex ? way1Tag_27 : _GEN_295; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_297 = 7'h1c == reqIndex ? way1Tag_28 : _GEN_296; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_298 = 7'h1d == reqIndex ? way1Tag_29 : _GEN_297; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_299 = 7'h1e == reqIndex ? way1Tag_30 : _GEN_298; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_300 = 7'h1f == reqIndex ? way1Tag_31 : _GEN_299; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_301 = 7'h20 == reqIndex ? way1Tag_32 : _GEN_300; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_302 = 7'h21 == reqIndex ? way1Tag_33 : _GEN_301; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_303 = 7'h22 == reqIndex ? way1Tag_34 : _GEN_302; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_304 = 7'h23 == reqIndex ? way1Tag_35 : _GEN_303; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_305 = 7'h24 == reqIndex ? way1Tag_36 : _GEN_304; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_306 = 7'h25 == reqIndex ? way1Tag_37 : _GEN_305; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_307 = 7'h26 == reqIndex ? way1Tag_38 : _GEN_306; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_308 = 7'h27 == reqIndex ? way1Tag_39 : _GEN_307; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_309 = 7'h28 == reqIndex ? way1Tag_40 : _GEN_308; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_310 = 7'h29 == reqIndex ? way1Tag_41 : _GEN_309; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_311 = 7'h2a == reqIndex ? way1Tag_42 : _GEN_310; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_312 = 7'h2b == reqIndex ? way1Tag_43 : _GEN_311; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_313 = 7'h2c == reqIndex ? way1Tag_44 : _GEN_312; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_314 = 7'h2d == reqIndex ? way1Tag_45 : _GEN_313; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_315 = 7'h2e == reqIndex ? way1Tag_46 : _GEN_314; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_316 = 7'h2f == reqIndex ? way1Tag_47 : _GEN_315; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_317 = 7'h30 == reqIndex ? way1Tag_48 : _GEN_316; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_318 = 7'h31 == reqIndex ? way1Tag_49 : _GEN_317; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_319 = 7'h32 == reqIndex ? way1Tag_50 : _GEN_318; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_320 = 7'h33 == reqIndex ? way1Tag_51 : _GEN_319; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_321 = 7'h34 == reqIndex ? way1Tag_52 : _GEN_320; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_322 = 7'h35 == reqIndex ? way1Tag_53 : _GEN_321; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_323 = 7'h36 == reqIndex ? way1Tag_54 : _GEN_322; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_324 = 7'h37 == reqIndex ? way1Tag_55 : _GEN_323; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_325 = 7'h38 == reqIndex ? way1Tag_56 : _GEN_324; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_326 = 7'h39 == reqIndex ? way1Tag_57 : _GEN_325; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_327 = 7'h3a == reqIndex ? way1Tag_58 : _GEN_326; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_328 = 7'h3b == reqIndex ? way1Tag_59 : _GEN_327; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_329 = 7'h3c == reqIndex ? way1Tag_60 : _GEN_328; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_330 = 7'h3d == reqIndex ? way1Tag_61 : _GEN_329; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_331 = 7'h3e == reqIndex ? way1Tag_62 : _GEN_330; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_332 = 7'h3f == reqIndex ? way1Tag_63 : _GEN_331; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_333 = 7'h40 == reqIndex ? way1Tag_64 : _GEN_332; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_334 = 7'h41 == reqIndex ? way1Tag_65 : _GEN_333; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_335 = 7'h42 == reqIndex ? way1Tag_66 : _GEN_334; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_336 = 7'h43 == reqIndex ? way1Tag_67 : _GEN_335; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_337 = 7'h44 == reqIndex ? way1Tag_68 : _GEN_336; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_338 = 7'h45 == reqIndex ? way1Tag_69 : _GEN_337; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_339 = 7'h46 == reqIndex ? way1Tag_70 : _GEN_338; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_340 = 7'h47 == reqIndex ? way1Tag_71 : _GEN_339; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_341 = 7'h48 == reqIndex ? way1Tag_72 : _GEN_340; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_342 = 7'h49 == reqIndex ? way1Tag_73 : _GEN_341; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_343 = 7'h4a == reqIndex ? way1Tag_74 : _GEN_342; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_344 = 7'h4b == reqIndex ? way1Tag_75 : _GEN_343; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_345 = 7'h4c == reqIndex ? way1Tag_76 : _GEN_344; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_346 = 7'h4d == reqIndex ? way1Tag_77 : _GEN_345; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_347 = 7'h4e == reqIndex ? way1Tag_78 : _GEN_346; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_348 = 7'h4f == reqIndex ? way1Tag_79 : _GEN_347; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_349 = 7'h50 == reqIndex ? way1Tag_80 : _GEN_348; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_350 = 7'h51 == reqIndex ? way1Tag_81 : _GEN_349; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_351 = 7'h52 == reqIndex ? way1Tag_82 : _GEN_350; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_352 = 7'h53 == reqIndex ? way1Tag_83 : _GEN_351; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_353 = 7'h54 == reqIndex ? way1Tag_84 : _GEN_352; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_354 = 7'h55 == reqIndex ? way1Tag_85 : _GEN_353; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_355 = 7'h56 == reqIndex ? way1Tag_86 : _GEN_354; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_356 = 7'h57 == reqIndex ? way1Tag_87 : _GEN_355; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_357 = 7'h58 == reqIndex ? way1Tag_88 : _GEN_356; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_358 = 7'h59 == reqIndex ? way1Tag_89 : _GEN_357; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_359 = 7'h5a == reqIndex ? way1Tag_90 : _GEN_358; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_360 = 7'h5b == reqIndex ? way1Tag_91 : _GEN_359; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_361 = 7'h5c == reqIndex ? way1Tag_92 : _GEN_360; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_362 = 7'h5d == reqIndex ? way1Tag_93 : _GEN_361; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_363 = 7'h5e == reqIndex ? way1Tag_94 : _GEN_362; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_364 = 7'h5f == reqIndex ? way1Tag_95 : _GEN_363; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_365 = 7'h60 == reqIndex ? way1Tag_96 : _GEN_364; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_366 = 7'h61 == reqIndex ? way1Tag_97 : _GEN_365; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_367 = 7'h62 == reqIndex ? way1Tag_98 : _GEN_366; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_368 = 7'h63 == reqIndex ? way1Tag_99 : _GEN_367; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_369 = 7'h64 == reqIndex ? way1Tag_100 : _GEN_368; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_370 = 7'h65 == reqIndex ? way1Tag_101 : _GEN_369; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_371 = 7'h66 == reqIndex ? way1Tag_102 : _GEN_370; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_372 = 7'h67 == reqIndex ? way1Tag_103 : _GEN_371; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_373 = 7'h68 == reqIndex ? way1Tag_104 : _GEN_372; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_374 = 7'h69 == reqIndex ? way1Tag_105 : _GEN_373; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_375 = 7'h6a == reqIndex ? way1Tag_106 : _GEN_374; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_376 = 7'h6b == reqIndex ? way1Tag_107 : _GEN_375; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_377 = 7'h6c == reqIndex ? way1Tag_108 : _GEN_376; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_378 = 7'h6d == reqIndex ? way1Tag_109 : _GEN_377; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_379 = 7'h6e == reqIndex ? way1Tag_110 : _GEN_378; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_380 = 7'h6f == reqIndex ? way1Tag_111 : _GEN_379; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_381 = 7'h70 == reqIndex ? way1Tag_112 : _GEN_380; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_382 = 7'h71 == reqIndex ? way1Tag_113 : _GEN_381; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_383 = 7'h72 == reqIndex ? way1Tag_114 : _GEN_382; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_384 = 7'h73 == reqIndex ? way1Tag_115 : _GEN_383; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_385 = 7'h74 == reqIndex ? way1Tag_116 : _GEN_384; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_386 = 7'h75 == reqIndex ? way1Tag_117 : _GEN_385; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_387 = 7'h76 == reqIndex ? way1Tag_118 : _GEN_386; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_388 = 7'h77 == reqIndex ? way1Tag_119 : _GEN_387; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_389 = 7'h78 == reqIndex ? way1Tag_120 : _GEN_388; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_390 = 7'h79 == reqIndex ? way1Tag_121 : _GEN_389; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_391 = 7'h7a == reqIndex ? way1Tag_122 : _GEN_390; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_392 = 7'h7b == reqIndex ? way1Tag_123 : _GEN_391; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_393 = 7'h7c == reqIndex ? way1Tag_124 : _GEN_392; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_394 = 7'h7d == reqIndex ? way1Tag_125 : _GEN_393; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_395 = 7'h7e == reqIndex ? way1Tag_126 : _GEN_394; // @[DCache.scala 125:{55,55}]
  wire [20:0] _GEN_396 = 7'h7f == reqIndex ? way1Tag_127 : _GEN_395; // @[DCache.scala 125:{55,55}]
  wire  way1Hit = _GEN_524 & _GEN_396 == reqTag; // @[DCache.scala 125:33]
  wire  cacheHitEn = way0Hit | way1Hit; // @[DCache.scala 126:26]
  wire  _cacheLineWay_T = way0Hit ? 1'h0 : 1'h1; // @[DCache.scala 132:38]
  wire  _ageWay0En_T = ~cacheHitEn; // @[DCache.scala 129:19]
  wire  _GEN_526 = 7'h1 == reqIndex ? way0Age_1 : way0Age_0; // @[DCache.scala 129:{53,53}]
  wire  _GEN_527 = 7'h2 == reqIndex ? way0Age_2 : _GEN_526; // @[DCache.scala 129:{53,53}]
  wire  _GEN_528 = 7'h3 == reqIndex ? way0Age_3 : _GEN_527; // @[DCache.scala 129:{53,53}]
  wire  _GEN_529 = 7'h4 == reqIndex ? way0Age_4 : _GEN_528; // @[DCache.scala 129:{53,53}]
  wire  _GEN_530 = 7'h5 == reqIndex ? way0Age_5 : _GEN_529; // @[DCache.scala 129:{53,53}]
  wire  _GEN_531 = 7'h6 == reqIndex ? way0Age_6 : _GEN_530; // @[DCache.scala 129:{53,53}]
  wire  _GEN_532 = 7'h7 == reqIndex ? way0Age_7 : _GEN_531; // @[DCache.scala 129:{53,53}]
  wire  _GEN_533 = 7'h8 == reqIndex ? way0Age_8 : _GEN_532; // @[DCache.scala 129:{53,53}]
  wire  _GEN_534 = 7'h9 == reqIndex ? way0Age_9 : _GEN_533; // @[DCache.scala 129:{53,53}]
  wire  _GEN_535 = 7'ha == reqIndex ? way0Age_10 : _GEN_534; // @[DCache.scala 129:{53,53}]
  wire  _GEN_536 = 7'hb == reqIndex ? way0Age_11 : _GEN_535; // @[DCache.scala 129:{53,53}]
  wire  _GEN_537 = 7'hc == reqIndex ? way0Age_12 : _GEN_536; // @[DCache.scala 129:{53,53}]
  wire  _GEN_538 = 7'hd == reqIndex ? way0Age_13 : _GEN_537; // @[DCache.scala 129:{53,53}]
  wire  _GEN_539 = 7'he == reqIndex ? way0Age_14 : _GEN_538; // @[DCache.scala 129:{53,53}]
  wire  _GEN_540 = 7'hf == reqIndex ? way0Age_15 : _GEN_539; // @[DCache.scala 129:{53,53}]
  wire  _GEN_541 = 7'h10 == reqIndex ? way0Age_16 : _GEN_540; // @[DCache.scala 129:{53,53}]
  wire  _GEN_542 = 7'h11 == reqIndex ? way0Age_17 : _GEN_541; // @[DCache.scala 129:{53,53}]
  wire  _GEN_543 = 7'h12 == reqIndex ? way0Age_18 : _GEN_542; // @[DCache.scala 129:{53,53}]
  wire  _GEN_544 = 7'h13 == reqIndex ? way0Age_19 : _GEN_543; // @[DCache.scala 129:{53,53}]
  wire  _GEN_545 = 7'h14 == reqIndex ? way0Age_20 : _GEN_544; // @[DCache.scala 129:{53,53}]
  wire  _GEN_546 = 7'h15 == reqIndex ? way0Age_21 : _GEN_545; // @[DCache.scala 129:{53,53}]
  wire  _GEN_547 = 7'h16 == reqIndex ? way0Age_22 : _GEN_546; // @[DCache.scala 129:{53,53}]
  wire  _GEN_548 = 7'h17 == reqIndex ? way0Age_23 : _GEN_547; // @[DCache.scala 129:{53,53}]
  wire  _GEN_549 = 7'h18 == reqIndex ? way0Age_24 : _GEN_548; // @[DCache.scala 129:{53,53}]
  wire  _GEN_550 = 7'h19 == reqIndex ? way0Age_25 : _GEN_549; // @[DCache.scala 129:{53,53}]
  wire  _GEN_551 = 7'h1a == reqIndex ? way0Age_26 : _GEN_550; // @[DCache.scala 129:{53,53}]
  wire  _GEN_552 = 7'h1b == reqIndex ? way0Age_27 : _GEN_551; // @[DCache.scala 129:{53,53}]
  wire  _GEN_553 = 7'h1c == reqIndex ? way0Age_28 : _GEN_552; // @[DCache.scala 129:{53,53}]
  wire  _GEN_554 = 7'h1d == reqIndex ? way0Age_29 : _GEN_553; // @[DCache.scala 129:{53,53}]
  wire  _GEN_555 = 7'h1e == reqIndex ? way0Age_30 : _GEN_554; // @[DCache.scala 129:{53,53}]
  wire  _GEN_556 = 7'h1f == reqIndex ? way0Age_31 : _GEN_555; // @[DCache.scala 129:{53,53}]
  wire  _GEN_557 = 7'h20 == reqIndex ? way0Age_32 : _GEN_556; // @[DCache.scala 129:{53,53}]
  wire  _GEN_558 = 7'h21 == reqIndex ? way0Age_33 : _GEN_557; // @[DCache.scala 129:{53,53}]
  wire  _GEN_559 = 7'h22 == reqIndex ? way0Age_34 : _GEN_558; // @[DCache.scala 129:{53,53}]
  wire  _GEN_560 = 7'h23 == reqIndex ? way0Age_35 : _GEN_559; // @[DCache.scala 129:{53,53}]
  wire  _GEN_561 = 7'h24 == reqIndex ? way0Age_36 : _GEN_560; // @[DCache.scala 129:{53,53}]
  wire  _GEN_562 = 7'h25 == reqIndex ? way0Age_37 : _GEN_561; // @[DCache.scala 129:{53,53}]
  wire  _GEN_563 = 7'h26 == reqIndex ? way0Age_38 : _GEN_562; // @[DCache.scala 129:{53,53}]
  wire  _GEN_564 = 7'h27 == reqIndex ? way0Age_39 : _GEN_563; // @[DCache.scala 129:{53,53}]
  wire  _GEN_565 = 7'h28 == reqIndex ? way0Age_40 : _GEN_564; // @[DCache.scala 129:{53,53}]
  wire  _GEN_566 = 7'h29 == reqIndex ? way0Age_41 : _GEN_565; // @[DCache.scala 129:{53,53}]
  wire  _GEN_567 = 7'h2a == reqIndex ? way0Age_42 : _GEN_566; // @[DCache.scala 129:{53,53}]
  wire  _GEN_568 = 7'h2b == reqIndex ? way0Age_43 : _GEN_567; // @[DCache.scala 129:{53,53}]
  wire  _GEN_569 = 7'h2c == reqIndex ? way0Age_44 : _GEN_568; // @[DCache.scala 129:{53,53}]
  wire  _GEN_570 = 7'h2d == reqIndex ? way0Age_45 : _GEN_569; // @[DCache.scala 129:{53,53}]
  wire  _GEN_571 = 7'h2e == reqIndex ? way0Age_46 : _GEN_570; // @[DCache.scala 129:{53,53}]
  wire  _GEN_572 = 7'h2f == reqIndex ? way0Age_47 : _GEN_571; // @[DCache.scala 129:{53,53}]
  wire  _GEN_573 = 7'h30 == reqIndex ? way0Age_48 : _GEN_572; // @[DCache.scala 129:{53,53}]
  wire  _GEN_574 = 7'h31 == reqIndex ? way0Age_49 : _GEN_573; // @[DCache.scala 129:{53,53}]
  wire  _GEN_575 = 7'h32 == reqIndex ? way0Age_50 : _GEN_574; // @[DCache.scala 129:{53,53}]
  wire  _GEN_576 = 7'h33 == reqIndex ? way0Age_51 : _GEN_575; // @[DCache.scala 129:{53,53}]
  wire  _GEN_577 = 7'h34 == reqIndex ? way0Age_52 : _GEN_576; // @[DCache.scala 129:{53,53}]
  wire  _GEN_578 = 7'h35 == reqIndex ? way0Age_53 : _GEN_577; // @[DCache.scala 129:{53,53}]
  wire  _GEN_579 = 7'h36 == reqIndex ? way0Age_54 : _GEN_578; // @[DCache.scala 129:{53,53}]
  wire  _GEN_580 = 7'h37 == reqIndex ? way0Age_55 : _GEN_579; // @[DCache.scala 129:{53,53}]
  wire  _GEN_581 = 7'h38 == reqIndex ? way0Age_56 : _GEN_580; // @[DCache.scala 129:{53,53}]
  wire  _GEN_582 = 7'h39 == reqIndex ? way0Age_57 : _GEN_581; // @[DCache.scala 129:{53,53}]
  wire  _GEN_583 = 7'h3a == reqIndex ? way0Age_58 : _GEN_582; // @[DCache.scala 129:{53,53}]
  wire  _GEN_584 = 7'h3b == reqIndex ? way0Age_59 : _GEN_583; // @[DCache.scala 129:{53,53}]
  wire  _GEN_585 = 7'h3c == reqIndex ? way0Age_60 : _GEN_584; // @[DCache.scala 129:{53,53}]
  wire  _GEN_586 = 7'h3d == reqIndex ? way0Age_61 : _GEN_585; // @[DCache.scala 129:{53,53}]
  wire  _GEN_587 = 7'h3e == reqIndex ? way0Age_62 : _GEN_586; // @[DCache.scala 129:{53,53}]
  wire  _GEN_588 = 7'h3f == reqIndex ? way0Age_63 : _GEN_587; // @[DCache.scala 129:{53,53}]
  wire  _GEN_589 = 7'h40 == reqIndex ? way0Age_64 : _GEN_588; // @[DCache.scala 129:{53,53}]
  wire  _GEN_590 = 7'h41 == reqIndex ? way0Age_65 : _GEN_589; // @[DCache.scala 129:{53,53}]
  wire  _GEN_591 = 7'h42 == reqIndex ? way0Age_66 : _GEN_590; // @[DCache.scala 129:{53,53}]
  wire  _GEN_592 = 7'h43 == reqIndex ? way0Age_67 : _GEN_591; // @[DCache.scala 129:{53,53}]
  wire  _GEN_593 = 7'h44 == reqIndex ? way0Age_68 : _GEN_592; // @[DCache.scala 129:{53,53}]
  wire  _GEN_594 = 7'h45 == reqIndex ? way0Age_69 : _GEN_593; // @[DCache.scala 129:{53,53}]
  wire  _GEN_595 = 7'h46 == reqIndex ? way0Age_70 : _GEN_594; // @[DCache.scala 129:{53,53}]
  wire  _GEN_596 = 7'h47 == reqIndex ? way0Age_71 : _GEN_595; // @[DCache.scala 129:{53,53}]
  wire  _GEN_597 = 7'h48 == reqIndex ? way0Age_72 : _GEN_596; // @[DCache.scala 129:{53,53}]
  wire  _GEN_598 = 7'h49 == reqIndex ? way0Age_73 : _GEN_597; // @[DCache.scala 129:{53,53}]
  wire  _GEN_599 = 7'h4a == reqIndex ? way0Age_74 : _GEN_598; // @[DCache.scala 129:{53,53}]
  wire  _GEN_600 = 7'h4b == reqIndex ? way0Age_75 : _GEN_599; // @[DCache.scala 129:{53,53}]
  wire  _GEN_601 = 7'h4c == reqIndex ? way0Age_76 : _GEN_600; // @[DCache.scala 129:{53,53}]
  wire  _GEN_602 = 7'h4d == reqIndex ? way0Age_77 : _GEN_601; // @[DCache.scala 129:{53,53}]
  wire  _GEN_603 = 7'h4e == reqIndex ? way0Age_78 : _GEN_602; // @[DCache.scala 129:{53,53}]
  wire  _GEN_604 = 7'h4f == reqIndex ? way0Age_79 : _GEN_603; // @[DCache.scala 129:{53,53}]
  wire  _GEN_605 = 7'h50 == reqIndex ? way0Age_80 : _GEN_604; // @[DCache.scala 129:{53,53}]
  wire  _GEN_606 = 7'h51 == reqIndex ? way0Age_81 : _GEN_605; // @[DCache.scala 129:{53,53}]
  wire  _GEN_607 = 7'h52 == reqIndex ? way0Age_82 : _GEN_606; // @[DCache.scala 129:{53,53}]
  wire  _GEN_608 = 7'h53 == reqIndex ? way0Age_83 : _GEN_607; // @[DCache.scala 129:{53,53}]
  wire  _GEN_609 = 7'h54 == reqIndex ? way0Age_84 : _GEN_608; // @[DCache.scala 129:{53,53}]
  wire  _GEN_610 = 7'h55 == reqIndex ? way0Age_85 : _GEN_609; // @[DCache.scala 129:{53,53}]
  wire  _GEN_611 = 7'h56 == reqIndex ? way0Age_86 : _GEN_610; // @[DCache.scala 129:{53,53}]
  wire  _GEN_612 = 7'h57 == reqIndex ? way0Age_87 : _GEN_611; // @[DCache.scala 129:{53,53}]
  wire  _GEN_613 = 7'h58 == reqIndex ? way0Age_88 : _GEN_612; // @[DCache.scala 129:{53,53}]
  wire  _GEN_614 = 7'h59 == reqIndex ? way0Age_89 : _GEN_613; // @[DCache.scala 129:{53,53}]
  wire  _GEN_615 = 7'h5a == reqIndex ? way0Age_90 : _GEN_614; // @[DCache.scala 129:{53,53}]
  wire  _GEN_616 = 7'h5b == reqIndex ? way0Age_91 : _GEN_615; // @[DCache.scala 129:{53,53}]
  wire  _GEN_617 = 7'h5c == reqIndex ? way0Age_92 : _GEN_616; // @[DCache.scala 129:{53,53}]
  wire  _GEN_618 = 7'h5d == reqIndex ? way0Age_93 : _GEN_617; // @[DCache.scala 129:{53,53}]
  wire  _GEN_619 = 7'h5e == reqIndex ? way0Age_94 : _GEN_618; // @[DCache.scala 129:{53,53}]
  wire  _GEN_620 = 7'h5f == reqIndex ? way0Age_95 : _GEN_619; // @[DCache.scala 129:{53,53}]
  wire  _GEN_621 = 7'h60 == reqIndex ? way0Age_96 : _GEN_620; // @[DCache.scala 129:{53,53}]
  wire  _GEN_622 = 7'h61 == reqIndex ? way0Age_97 : _GEN_621; // @[DCache.scala 129:{53,53}]
  wire  _GEN_623 = 7'h62 == reqIndex ? way0Age_98 : _GEN_622; // @[DCache.scala 129:{53,53}]
  wire  _GEN_624 = 7'h63 == reqIndex ? way0Age_99 : _GEN_623; // @[DCache.scala 129:{53,53}]
  wire  _GEN_625 = 7'h64 == reqIndex ? way0Age_100 : _GEN_624; // @[DCache.scala 129:{53,53}]
  wire  _GEN_626 = 7'h65 == reqIndex ? way0Age_101 : _GEN_625; // @[DCache.scala 129:{53,53}]
  wire  _GEN_627 = 7'h66 == reqIndex ? way0Age_102 : _GEN_626; // @[DCache.scala 129:{53,53}]
  wire  _GEN_628 = 7'h67 == reqIndex ? way0Age_103 : _GEN_627; // @[DCache.scala 129:{53,53}]
  wire  _GEN_629 = 7'h68 == reqIndex ? way0Age_104 : _GEN_628; // @[DCache.scala 129:{53,53}]
  wire  _GEN_630 = 7'h69 == reqIndex ? way0Age_105 : _GEN_629; // @[DCache.scala 129:{53,53}]
  wire  _GEN_631 = 7'h6a == reqIndex ? way0Age_106 : _GEN_630; // @[DCache.scala 129:{53,53}]
  wire  _GEN_632 = 7'h6b == reqIndex ? way0Age_107 : _GEN_631; // @[DCache.scala 129:{53,53}]
  wire  _GEN_633 = 7'h6c == reqIndex ? way0Age_108 : _GEN_632; // @[DCache.scala 129:{53,53}]
  wire  _GEN_634 = 7'h6d == reqIndex ? way0Age_109 : _GEN_633; // @[DCache.scala 129:{53,53}]
  wire  _GEN_635 = 7'h6e == reqIndex ? way0Age_110 : _GEN_634; // @[DCache.scala 129:{53,53}]
  wire  _GEN_636 = 7'h6f == reqIndex ? way0Age_111 : _GEN_635; // @[DCache.scala 129:{53,53}]
  wire  _GEN_637 = 7'h70 == reqIndex ? way0Age_112 : _GEN_636; // @[DCache.scala 129:{53,53}]
  wire  _GEN_638 = 7'h71 == reqIndex ? way0Age_113 : _GEN_637; // @[DCache.scala 129:{53,53}]
  wire  _GEN_639 = 7'h72 == reqIndex ? way0Age_114 : _GEN_638; // @[DCache.scala 129:{53,53}]
  wire  _GEN_640 = 7'h73 == reqIndex ? way0Age_115 : _GEN_639; // @[DCache.scala 129:{53,53}]
  wire  _GEN_641 = 7'h74 == reqIndex ? way0Age_116 : _GEN_640; // @[DCache.scala 129:{53,53}]
  wire  _GEN_642 = 7'h75 == reqIndex ? way0Age_117 : _GEN_641; // @[DCache.scala 129:{53,53}]
  wire  _GEN_643 = 7'h76 == reqIndex ? way0Age_118 : _GEN_642; // @[DCache.scala 129:{53,53}]
  wire  _GEN_644 = 7'h77 == reqIndex ? way0Age_119 : _GEN_643; // @[DCache.scala 129:{53,53}]
  wire  _GEN_645 = 7'h78 == reqIndex ? way0Age_120 : _GEN_644; // @[DCache.scala 129:{53,53}]
  wire  _GEN_646 = 7'h79 == reqIndex ? way0Age_121 : _GEN_645; // @[DCache.scala 129:{53,53}]
  wire  _GEN_647 = 7'h7a == reqIndex ? way0Age_122 : _GEN_646; // @[DCache.scala 129:{53,53}]
  wire  _GEN_648 = 7'h7b == reqIndex ? way0Age_123 : _GEN_647; // @[DCache.scala 129:{53,53}]
  wire  _GEN_649 = 7'h7c == reqIndex ? way0Age_124 : _GEN_648; // @[DCache.scala 129:{53,53}]
  wire  _GEN_650 = 7'h7d == reqIndex ? way0Age_125 : _GEN_649; // @[DCache.scala 129:{53,53}]
  wire  _GEN_651 = 7'h7e == reqIndex ? way0Age_126 : _GEN_650; // @[DCache.scala 129:{53,53}]
  wire  _GEN_652 = 7'h7f == reqIndex ? way0Age_127 : _GEN_651; // @[DCache.scala 129:{53,53}]
  wire  ageWay0En = ~cacheHitEn & ~_GEN_652; // @[DCache.scala 129:31]
  wire  _cacheLineWay_T_1 = ageWay0En ? 1'h0 : 1'h1; // @[DCache.scala 132:62]
  wire  cacheLineWay = cacheHitEn ? _cacheLineWay_T : _cacheLineWay_T_1; // @[DCache.scala 132:22]
  wire  _cacheDirtyEn_T = ~cacheLineWay; // @[DCache.scala 136:36]
  wire  _GEN_782 = 7'h1 == reqIndex ? way0Dirty_1 : way0Dirty_0; // @[DCache.scala 136:{22,22}]
  wire  _GEN_783 = 7'h2 == reqIndex ? way0Dirty_2 : _GEN_782; // @[DCache.scala 136:{22,22}]
  wire  _GEN_784 = 7'h3 == reqIndex ? way0Dirty_3 : _GEN_783; // @[DCache.scala 136:{22,22}]
  wire  _GEN_785 = 7'h4 == reqIndex ? way0Dirty_4 : _GEN_784; // @[DCache.scala 136:{22,22}]
  wire  _GEN_786 = 7'h5 == reqIndex ? way0Dirty_5 : _GEN_785; // @[DCache.scala 136:{22,22}]
  wire  _GEN_787 = 7'h6 == reqIndex ? way0Dirty_6 : _GEN_786; // @[DCache.scala 136:{22,22}]
  wire  _GEN_788 = 7'h7 == reqIndex ? way0Dirty_7 : _GEN_787; // @[DCache.scala 136:{22,22}]
  wire  _GEN_789 = 7'h8 == reqIndex ? way0Dirty_8 : _GEN_788; // @[DCache.scala 136:{22,22}]
  wire  _GEN_790 = 7'h9 == reqIndex ? way0Dirty_9 : _GEN_789; // @[DCache.scala 136:{22,22}]
  wire  _GEN_791 = 7'ha == reqIndex ? way0Dirty_10 : _GEN_790; // @[DCache.scala 136:{22,22}]
  wire  _GEN_792 = 7'hb == reqIndex ? way0Dirty_11 : _GEN_791; // @[DCache.scala 136:{22,22}]
  wire  _GEN_793 = 7'hc == reqIndex ? way0Dirty_12 : _GEN_792; // @[DCache.scala 136:{22,22}]
  wire  _GEN_794 = 7'hd == reqIndex ? way0Dirty_13 : _GEN_793; // @[DCache.scala 136:{22,22}]
  wire  _GEN_795 = 7'he == reqIndex ? way0Dirty_14 : _GEN_794; // @[DCache.scala 136:{22,22}]
  wire  _GEN_796 = 7'hf == reqIndex ? way0Dirty_15 : _GEN_795; // @[DCache.scala 136:{22,22}]
  wire  _GEN_797 = 7'h10 == reqIndex ? way0Dirty_16 : _GEN_796; // @[DCache.scala 136:{22,22}]
  wire  _GEN_798 = 7'h11 == reqIndex ? way0Dirty_17 : _GEN_797; // @[DCache.scala 136:{22,22}]
  wire  _GEN_799 = 7'h12 == reqIndex ? way0Dirty_18 : _GEN_798; // @[DCache.scala 136:{22,22}]
  wire  _GEN_800 = 7'h13 == reqIndex ? way0Dirty_19 : _GEN_799; // @[DCache.scala 136:{22,22}]
  wire  _GEN_801 = 7'h14 == reqIndex ? way0Dirty_20 : _GEN_800; // @[DCache.scala 136:{22,22}]
  wire  _GEN_802 = 7'h15 == reqIndex ? way0Dirty_21 : _GEN_801; // @[DCache.scala 136:{22,22}]
  wire  _GEN_803 = 7'h16 == reqIndex ? way0Dirty_22 : _GEN_802; // @[DCache.scala 136:{22,22}]
  wire  _GEN_804 = 7'h17 == reqIndex ? way0Dirty_23 : _GEN_803; // @[DCache.scala 136:{22,22}]
  wire  _GEN_805 = 7'h18 == reqIndex ? way0Dirty_24 : _GEN_804; // @[DCache.scala 136:{22,22}]
  wire  _GEN_806 = 7'h19 == reqIndex ? way0Dirty_25 : _GEN_805; // @[DCache.scala 136:{22,22}]
  wire  _GEN_807 = 7'h1a == reqIndex ? way0Dirty_26 : _GEN_806; // @[DCache.scala 136:{22,22}]
  wire  _GEN_808 = 7'h1b == reqIndex ? way0Dirty_27 : _GEN_807; // @[DCache.scala 136:{22,22}]
  wire  _GEN_809 = 7'h1c == reqIndex ? way0Dirty_28 : _GEN_808; // @[DCache.scala 136:{22,22}]
  wire  _GEN_810 = 7'h1d == reqIndex ? way0Dirty_29 : _GEN_809; // @[DCache.scala 136:{22,22}]
  wire  _GEN_811 = 7'h1e == reqIndex ? way0Dirty_30 : _GEN_810; // @[DCache.scala 136:{22,22}]
  wire  _GEN_812 = 7'h1f == reqIndex ? way0Dirty_31 : _GEN_811; // @[DCache.scala 136:{22,22}]
  wire  _GEN_813 = 7'h20 == reqIndex ? way0Dirty_32 : _GEN_812; // @[DCache.scala 136:{22,22}]
  wire  _GEN_814 = 7'h21 == reqIndex ? way0Dirty_33 : _GEN_813; // @[DCache.scala 136:{22,22}]
  wire  _GEN_815 = 7'h22 == reqIndex ? way0Dirty_34 : _GEN_814; // @[DCache.scala 136:{22,22}]
  wire  _GEN_816 = 7'h23 == reqIndex ? way0Dirty_35 : _GEN_815; // @[DCache.scala 136:{22,22}]
  wire  _GEN_817 = 7'h24 == reqIndex ? way0Dirty_36 : _GEN_816; // @[DCache.scala 136:{22,22}]
  wire  _GEN_818 = 7'h25 == reqIndex ? way0Dirty_37 : _GEN_817; // @[DCache.scala 136:{22,22}]
  wire  _GEN_819 = 7'h26 == reqIndex ? way0Dirty_38 : _GEN_818; // @[DCache.scala 136:{22,22}]
  wire  _GEN_820 = 7'h27 == reqIndex ? way0Dirty_39 : _GEN_819; // @[DCache.scala 136:{22,22}]
  wire  _GEN_821 = 7'h28 == reqIndex ? way0Dirty_40 : _GEN_820; // @[DCache.scala 136:{22,22}]
  wire  _GEN_822 = 7'h29 == reqIndex ? way0Dirty_41 : _GEN_821; // @[DCache.scala 136:{22,22}]
  wire  _GEN_823 = 7'h2a == reqIndex ? way0Dirty_42 : _GEN_822; // @[DCache.scala 136:{22,22}]
  wire  _GEN_824 = 7'h2b == reqIndex ? way0Dirty_43 : _GEN_823; // @[DCache.scala 136:{22,22}]
  wire  _GEN_825 = 7'h2c == reqIndex ? way0Dirty_44 : _GEN_824; // @[DCache.scala 136:{22,22}]
  wire  _GEN_826 = 7'h2d == reqIndex ? way0Dirty_45 : _GEN_825; // @[DCache.scala 136:{22,22}]
  wire  _GEN_827 = 7'h2e == reqIndex ? way0Dirty_46 : _GEN_826; // @[DCache.scala 136:{22,22}]
  wire  _GEN_828 = 7'h2f == reqIndex ? way0Dirty_47 : _GEN_827; // @[DCache.scala 136:{22,22}]
  wire  _GEN_829 = 7'h30 == reqIndex ? way0Dirty_48 : _GEN_828; // @[DCache.scala 136:{22,22}]
  wire  _GEN_830 = 7'h31 == reqIndex ? way0Dirty_49 : _GEN_829; // @[DCache.scala 136:{22,22}]
  wire  _GEN_831 = 7'h32 == reqIndex ? way0Dirty_50 : _GEN_830; // @[DCache.scala 136:{22,22}]
  wire  _GEN_832 = 7'h33 == reqIndex ? way0Dirty_51 : _GEN_831; // @[DCache.scala 136:{22,22}]
  wire  _GEN_833 = 7'h34 == reqIndex ? way0Dirty_52 : _GEN_832; // @[DCache.scala 136:{22,22}]
  wire  _GEN_834 = 7'h35 == reqIndex ? way0Dirty_53 : _GEN_833; // @[DCache.scala 136:{22,22}]
  wire  _GEN_835 = 7'h36 == reqIndex ? way0Dirty_54 : _GEN_834; // @[DCache.scala 136:{22,22}]
  wire  _GEN_836 = 7'h37 == reqIndex ? way0Dirty_55 : _GEN_835; // @[DCache.scala 136:{22,22}]
  wire  _GEN_837 = 7'h38 == reqIndex ? way0Dirty_56 : _GEN_836; // @[DCache.scala 136:{22,22}]
  wire  _GEN_838 = 7'h39 == reqIndex ? way0Dirty_57 : _GEN_837; // @[DCache.scala 136:{22,22}]
  wire  _GEN_839 = 7'h3a == reqIndex ? way0Dirty_58 : _GEN_838; // @[DCache.scala 136:{22,22}]
  wire  _GEN_840 = 7'h3b == reqIndex ? way0Dirty_59 : _GEN_839; // @[DCache.scala 136:{22,22}]
  wire  _GEN_841 = 7'h3c == reqIndex ? way0Dirty_60 : _GEN_840; // @[DCache.scala 136:{22,22}]
  wire  _GEN_842 = 7'h3d == reqIndex ? way0Dirty_61 : _GEN_841; // @[DCache.scala 136:{22,22}]
  wire  _GEN_843 = 7'h3e == reqIndex ? way0Dirty_62 : _GEN_842; // @[DCache.scala 136:{22,22}]
  wire  _GEN_844 = 7'h3f == reqIndex ? way0Dirty_63 : _GEN_843; // @[DCache.scala 136:{22,22}]
  wire  _GEN_845 = 7'h40 == reqIndex ? way0Dirty_64 : _GEN_844; // @[DCache.scala 136:{22,22}]
  wire  _GEN_846 = 7'h41 == reqIndex ? way0Dirty_65 : _GEN_845; // @[DCache.scala 136:{22,22}]
  wire  _GEN_847 = 7'h42 == reqIndex ? way0Dirty_66 : _GEN_846; // @[DCache.scala 136:{22,22}]
  wire  _GEN_848 = 7'h43 == reqIndex ? way0Dirty_67 : _GEN_847; // @[DCache.scala 136:{22,22}]
  wire  _GEN_849 = 7'h44 == reqIndex ? way0Dirty_68 : _GEN_848; // @[DCache.scala 136:{22,22}]
  wire  _GEN_850 = 7'h45 == reqIndex ? way0Dirty_69 : _GEN_849; // @[DCache.scala 136:{22,22}]
  wire  _GEN_851 = 7'h46 == reqIndex ? way0Dirty_70 : _GEN_850; // @[DCache.scala 136:{22,22}]
  wire  _GEN_852 = 7'h47 == reqIndex ? way0Dirty_71 : _GEN_851; // @[DCache.scala 136:{22,22}]
  wire  _GEN_853 = 7'h48 == reqIndex ? way0Dirty_72 : _GEN_852; // @[DCache.scala 136:{22,22}]
  wire  _GEN_854 = 7'h49 == reqIndex ? way0Dirty_73 : _GEN_853; // @[DCache.scala 136:{22,22}]
  wire  _GEN_855 = 7'h4a == reqIndex ? way0Dirty_74 : _GEN_854; // @[DCache.scala 136:{22,22}]
  wire  _GEN_856 = 7'h4b == reqIndex ? way0Dirty_75 : _GEN_855; // @[DCache.scala 136:{22,22}]
  wire  _GEN_857 = 7'h4c == reqIndex ? way0Dirty_76 : _GEN_856; // @[DCache.scala 136:{22,22}]
  wire  _GEN_858 = 7'h4d == reqIndex ? way0Dirty_77 : _GEN_857; // @[DCache.scala 136:{22,22}]
  wire  _GEN_859 = 7'h4e == reqIndex ? way0Dirty_78 : _GEN_858; // @[DCache.scala 136:{22,22}]
  wire  _GEN_860 = 7'h4f == reqIndex ? way0Dirty_79 : _GEN_859; // @[DCache.scala 136:{22,22}]
  wire  _GEN_861 = 7'h50 == reqIndex ? way0Dirty_80 : _GEN_860; // @[DCache.scala 136:{22,22}]
  wire  _GEN_862 = 7'h51 == reqIndex ? way0Dirty_81 : _GEN_861; // @[DCache.scala 136:{22,22}]
  wire  _GEN_863 = 7'h52 == reqIndex ? way0Dirty_82 : _GEN_862; // @[DCache.scala 136:{22,22}]
  wire  _GEN_864 = 7'h53 == reqIndex ? way0Dirty_83 : _GEN_863; // @[DCache.scala 136:{22,22}]
  wire  _GEN_865 = 7'h54 == reqIndex ? way0Dirty_84 : _GEN_864; // @[DCache.scala 136:{22,22}]
  wire  _GEN_866 = 7'h55 == reqIndex ? way0Dirty_85 : _GEN_865; // @[DCache.scala 136:{22,22}]
  wire  _GEN_867 = 7'h56 == reqIndex ? way0Dirty_86 : _GEN_866; // @[DCache.scala 136:{22,22}]
  wire  _GEN_868 = 7'h57 == reqIndex ? way0Dirty_87 : _GEN_867; // @[DCache.scala 136:{22,22}]
  wire  _GEN_869 = 7'h58 == reqIndex ? way0Dirty_88 : _GEN_868; // @[DCache.scala 136:{22,22}]
  wire  _GEN_870 = 7'h59 == reqIndex ? way0Dirty_89 : _GEN_869; // @[DCache.scala 136:{22,22}]
  wire  _GEN_871 = 7'h5a == reqIndex ? way0Dirty_90 : _GEN_870; // @[DCache.scala 136:{22,22}]
  wire  _GEN_872 = 7'h5b == reqIndex ? way0Dirty_91 : _GEN_871; // @[DCache.scala 136:{22,22}]
  wire  _GEN_873 = 7'h5c == reqIndex ? way0Dirty_92 : _GEN_872; // @[DCache.scala 136:{22,22}]
  wire  _GEN_874 = 7'h5d == reqIndex ? way0Dirty_93 : _GEN_873; // @[DCache.scala 136:{22,22}]
  wire  _GEN_875 = 7'h5e == reqIndex ? way0Dirty_94 : _GEN_874; // @[DCache.scala 136:{22,22}]
  wire  _GEN_876 = 7'h5f == reqIndex ? way0Dirty_95 : _GEN_875; // @[DCache.scala 136:{22,22}]
  wire  _GEN_877 = 7'h60 == reqIndex ? way0Dirty_96 : _GEN_876; // @[DCache.scala 136:{22,22}]
  wire  _GEN_878 = 7'h61 == reqIndex ? way0Dirty_97 : _GEN_877; // @[DCache.scala 136:{22,22}]
  wire  _GEN_879 = 7'h62 == reqIndex ? way0Dirty_98 : _GEN_878; // @[DCache.scala 136:{22,22}]
  wire  _GEN_880 = 7'h63 == reqIndex ? way0Dirty_99 : _GEN_879; // @[DCache.scala 136:{22,22}]
  wire  _GEN_881 = 7'h64 == reqIndex ? way0Dirty_100 : _GEN_880; // @[DCache.scala 136:{22,22}]
  wire  _GEN_882 = 7'h65 == reqIndex ? way0Dirty_101 : _GEN_881; // @[DCache.scala 136:{22,22}]
  wire  _GEN_883 = 7'h66 == reqIndex ? way0Dirty_102 : _GEN_882; // @[DCache.scala 136:{22,22}]
  wire  _GEN_884 = 7'h67 == reqIndex ? way0Dirty_103 : _GEN_883; // @[DCache.scala 136:{22,22}]
  wire  _GEN_885 = 7'h68 == reqIndex ? way0Dirty_104 : _GEN_884; // @[DCache.scala 136:{22,22}]
  wire  _GEN_886 = 7'h69 == reqIndex ? way0Dirty_105 : _GEN_885; // @[DCache.scala 136:{22,22}]
  wire  _GEN_887 = 7'h6a == reqIndex ? way0Dirty_106 : _GEN_886; // @[DCache.scala 136:{22,22}]
  wire  _GEN_888 = 7'h6b == reqIndex ? way0Dirty_107 : _GEN_887; // @[DCache.scala 136:{22,22}]
  wire  _GEN_889 = 7'h6c == reqIndex ? way0Dirty_108 : _GEN_888; // @[DCache.scala 136:{22,22}]
  wire  _GEN_890 = 7'h6d == reqIndex ? way0Dirty_109 : _GEN_889; // @[DCache.scala 136:{22,22}]
  wire  _GEN_891 = 7'h6e == reqIndex ? way0Dirty_110 : _GEN_890; // @[DCache.scala 136:{22,22}]
  wire  _GEN_892 = 7'h6f == reqIndex ? way0Dirty_111 : _GEN_891; // @[DCache.scala 136:{22,22}]
  wire  _GEN_893 = 7'h70 == reqIndex ? way0Dirty_112 : _GEN_892; // @[DCache.scala 136:{22,22}]
  wire  _GEN_894 = 7'h71 == reqIndex ? way0Dirty_113 : _GEN_893; // @[DCache.scala 136:{22,22}]
  wire  _GEN_895 = 7'h72 == reqIndex ? way0Dirty_114 : _GEN_894; // @[DCache.scala 136:{22,22}]
  wire  _GEN_896 = 7'h73 == reqIndex ? way0Dirty_115 : _GEN_895; // @[DCache.scala 136:{22,22}]
  wire  _GEN_897 = 7'h74 == reqIndex ? way0Dirty_116 : _GEN_896; // @[DCache.scala 136:{22,22}]
  wire  _GEN_898 = 7'h75 == reqIndex ? way0Dirty_117 : _GEN_897; // @[DCache.scala 136:{22,22}]
  wire  _GEN_899 = 7'h76 == reqIndex ? way0Dirty_118 : _GEN_898; // @[DCache.scala 136:{22,22}]
  wire  _GEN_900 = 7'h77 == reqIndex ? way0Dirty_119 : _GEN_899; // @[DCache.scala 136:{22,22}]
  wire  _GEN_901 = 7'h78 == reqIndex ? way0Dirty_120 : _GEN_900; // @[DCache.scala 136:{22,22}]
  wire  _GEN_902 = 7'h79 == reqIndex ? way0Dirty_121 : _GEN_901; // @[DCache.scala 136:{22,22}]
  wire  _GEN_903 = 7'h7a == reqIndex ? way0Dirty_122 : _GEN_902; // @[DCache.scala 136:{22,22}]
  wire  _GEN_904 = 7'h7b == reqIndex ? way0Dirty_123 : _GEN_903; // @[DCache.scala 136:{22,22}]
  wire  _GEN_905 = 7'h7c == reqIndex ? way0Dirty_124 : _GEN_904; // @[DCache.scala 136:{22,22}]
  wire  _GEN_906 = 7'h7d == reqIndex ? way0Dirty_125 : _GEN_905; // @[DCache.scala 136:{22,22}]
  wire  _GEN_907 = 7'h7e == reqIndex ? way0Dirty_126 : _GEN_906; // @[DCache.scala 136:{22,22}]
  wire  _GEN_908 = 7'h7f == reqIndex ? way0Dirty_127 : _GEN_907; // @[DCache.scala 136:{22,22}]
  wire  _GEN_910 = 7'h1 == reqIndex ? way1Dirty_1 : way1Dirty_0; // @[DCache.scala 136:{22,22}]
  wire  _GEN_911 = 7'h2 == reqIndex ? way1Dirty_2 : _GEN_910; // @[DCache.scala 136:{22,22}]
  wire  _GEN_912 = 7'h3 == reqIndex ? way1Dirty_3 : _GEN_911; // @[DCache.scala 136:{22,22}]
  wire  _GEN_913 = 7'h4 == reqIndex ? way1Dirty_4 : _GEN_912; // @[DCache.scala 136:{22,22}]
  wire  _GEN_914 = 7'h5 == reqIndex ? way1Dirty_5 : _GEN_913; // @[DCache.scala 136:{22,22}]
  wire  _GEN_915 = 7'h6 == reqIndex ? way1Dirty_6 : _GEN_914; // @[DCache.scala 136:{22,22}]
  wire  _GEN_916 = 7'h7 == reqIndex ? way1Dirty_7 : _GEN_915; // @[DCache.scala 136:{22,22}]
  wire  _GEN_917 = 7'h8 == reqIndex ? way1Dirty_8 : _GEN_916; // @[DCache.scala 136:{22,22}]
  wire  _GEN_918 = 7'h9 == reqIndex ? way1Dirty_9 : _GEN_917; // @[DCache.scala 136:{22,22}]
  wire  _GEN_919 = 7'ha == reqIndex ? way1Dirty_10 : _GEN_918; // @[DCache.scala 136:{22,22}]
  wire  _GEN_920 = 7'hb == reqIndex ? way1Dirty_11 : _GEN_919; // @[DCache.scala 136:{22,22}]
  wire  _GEN_921 = 7'hc == reqIndex ? way1Dirty_12 : _GEN_920; // @[DCache.scala 136:{22,22}]
  wire  _GEN_922 = 7'hd == reqIndex ? way1Dirty_13 : _GEN_921; // @[DCache.scala 136:{22,22}]
  wire  _GEN_923 = 7'he == reqIndex ? way1Dirty_14 : _GEN_922; // @[DCache.scala 136:{22,22}]
  wire  _GEN_924 = 7'hf == reqIndex ? way1Dirty_15 : _GEN_923; // @[DCache.scala 136:{22,22}]
  wire  _GEN_925 = 7'h10 == reqIndex ? way1Dirty_16 : _GEN_924; // @[DCache.scala 136:{22,22}]
  wire  _GEN_926 = 7'h11 == reqIndex ? way1Dirty_17 : _GEN_925; // @[DCache.scala 136:{22,22}]
  wire  _GEN_927 = 7'h12 == reqIndex ? way1Dirty_18 : _GEN_926; // @[DCache.scala 136:{22,22}]
  wire  _GEN_928 = 7'h13 == reqIndex ? way1Dirty_19 : _GEN_927; // @[DCache.scala 136:{22,22}]
  wire  _GEN_929 = 7'h14 == reqIndex ? way1Dirty_20 : _GEN_928; // @[DCache.scala 136:{22,22}]
  wire  _GEN_930 = 7'h15 == reqIndex ? way1Dirty_21 : _GEN_929; // @[DCache.scala 136:{22,22}]
  wire  _GEN_931 = 7'h16 == reqIndex ? way1Dirty_22 : _GEN_930; // @[DCache.scala 136:{22,22}]
  wire  _GEN_932 = 7'h17 == reqIndex ? way1Dirty_23 : _GEN_931; // @[DCache.scala 136:{22,22}]
  wire  _GEN_933 = 7'h18 == reqIndex ? way1Dirty_24 : _GEN_932; // @[DCache.scala 136:{22,22}]
  wire  _GEN_934 = 7'h19 == reqIndex ? way1Dirty_25 : _GEN_933; // @[DCache.scala 136:{22,22}]
  wire  _GEN_935 = 7'h1a == reqIndex ? way1Dirty_26 : _GEN_934; // @[DCache.scala 136:{22,22}]
  wire  _GEN_936 = 7'h1b == reqIndex ? way1Dirty_27 : _GEN_935; // @[DCache.scala 136:{22,22}]
  wire  _GEN_937 = 7'h1c == reqIndex ? way1Dirty_28 : _GEN_936; // @[DCache.scala 136:{22,22}]
  wire  _GEN_938 = 7'h1d == reqIndex ? way1Dirty_29 : _GEN_937; // @[DCache.scala 136:{22,22}]
  wire  _GEN_939 = 7'h1e == reqIndex ? way1Dirty_30 : _GEN_938; // @[DCache.scala 136:{22,22}]
  wire  _GEN_940 = 7'h1f == reqIndex ? way1Dirty_31 : _GEN_939; // @[DCache.scala 136:{22,22}]
  wire  _GEN_941 = 7'h20 == reqIndex ? way1Dirty_32 : _GEN_940; // @[DCache.scala 136:{22,22}]
  wire  _GEN_942 = 7'h21 == reqIndex ? way1Dirty_33 : _GEN_941; // @[DCache.scala 136:{22,22}]
  wire  _GEN_943 = 7'h22 == reqIndex ? way1Dirty_34 : _GEN_942; // @[DCache.scala 136:{22,22}]
  wire  _GEN_944 = 7'h23 == reqIndex ? way1Dirty_35 : _GEN_943; // @[DCache.scala 136:{22,22}]
  wire  _GEN_945 = 7'h24 == reqIndex ? way1Dirty_36 : _GEN_944; // @[DCache.scala 136:{22,22}]
  wire  _GEN_946 = 7'h25 == reqIndex ? way1Dirty_37 : _GEN_945; // @[DCache.scala 136:{22,22}]
  wire  _GEN_947 = 7'h26 == reqIndex ? way1Dirty_38 : _GEN_946; // @[DCache.scala 136:{22,22}]
  wire  _GEN_948 = 7'h27 == reqIndex ? way1Dirty_39 : _GEN_947; // @[DCache.scala 136:{22,22}]
  wire  _GEN_949 = 7'h28 == reqIndex ? way1Dirty_40 : _GEN_948; // @[DCache.scala 136:{22,22}]
  wire  _GEN_950 = 7'h29 == reqIndex ? way1Dirty_41 : _GEN_949; // @[DCache.scala 136:{22,22}]
  wire  _GEN_951 = 7'h2a == reqIndex ? way1Dirty_42 : _GEN_950; // @[DCache.scala 136:{22,22}]
  wire  _GEN_952 = 7'h2b == reqIndex ? way1Dirty_43 : _GEN_951; // @[DCache.scala 136:{22,22}]
  wire  _GEN_953 = 7'h2c == reqIndex ? way1Dirty_44 : _GEN_952; // @[DCache.scala 136:{22,22}]
  wire  _GEN_954 = 7'h2d == reqIndex ? way1Dirty_45 : _GEN_953; // @[DCache.scala 136:{22,22}]
  wire  _GEN_955 = 7'h2e == reqIndex ? way1Dirty_46 : _GEN_954; // @[DCache.scala 136:{22,22}]
  wire  _GEN_956 = 7'h2f == reqIndex ? way1Dirty_47 : _GEN_955; // @[DCache.scala 136:{22,22}]
  wire  _GEN_957 = 7'h30 == reqIndex ? way1Dirty_48 : _GEN_956; // @[DCache.scala 136:{22,22}]
  wire  _GEN_958 = 7'h31 == reqIndex ? way1Dirty_49 : _GEN_957; // @[DCache.scala 136:{22,22}]
  wire  _GEN_959 = 7'h32 == reqIndex ? way1Dirty_50 : _GEN_958; // @[DCache.scala 136:{22,22}]
  wire  _GEN_960 = 7'h33 == reqIndex ? way1Dirty_51 : _GEN_959; // @[DCache.scala 136:{22,22}]
  wire  _GEN_961 = 7'h34 == reqIndex ? way1Dirty_52 : _GEN_960; // @[DCache.scala 136:{22,22}]
  wire  _GEN_962 = 7'h35 == reqIndex ? way1Dirty_53 : _GEN_961; // @[DCache.scala 136:{22,22}]
  wire  _GEN_963 = 7'h36 == reqIndex ? way1Dirty_54 : _GEN_962; // @[DCache.scala 136:{22,22}]
  wire  _GEN_964 = 7'h37 == reqIndex ? way1Dirty_55 : _GEN_963; // @[DCache.scala 136:{22,22}]
  wire  _GEN_965 = 7'h38 == reqIndex ? way1Dirty_56 : _GEN_964; // @[DCache.scala 136:{22,22}]
  wire  _GEN_966 = 7'h39 == reqIndex ? way1Dirty_57 : _GEN_965; // @[DCache.scala 136:{22,22}]
  wire  _GEN_967 = 7'h3a == reqIndex ? way1Dirty_58 : _GEN_966; // @[DCache.scala 136:{22,22}]
  wire  _GEN_968 = 7'h3b == reqIndex ? way1Dirty_59 : _GEN_967; // @[DCache.scala 136:{22,22}]
  wire  _GEN_969 = 7'h3c == reqIndex ? way1Dirty_60 : _GEN_968; // @[DCache.scala 136:{22,22}]
  wire  _GEN_970 = 7'h3d == reqIndex ? way1Dirty_61 : _GEN_969; // @[DCache.scala 136:{22,22}]
  wire  _GEN_971 = 7'h3e == reqIndex ? way1Dirty_62 : _GEN_970; // @[DCache.scala 136:{22,22}]
  wire  _GEN_972 = 7'h3f == reqIndex ? way1Dirty_63 : _GEN_971; // @[DCache.scala 136:{22,22}]
  wire  _GEN_973 = 7'h40 == reqIndex ? way1Dirty_64 : _GEN_972; // @[DCache.scala 136:{22,22}]
  wire  _GEN_974 = 7'h41 == reqIndex ? way1Dirty_65 : _GEN_973; // @[DCache.scala 136:{22,22}]
  wire  _GEN_975 = 7'h42 == reqIndex ? way1Dirty_66 : _GEN_974; // @[DCache.scala 136:{22,22}]
  wire  _GEN_976 = 7'h43 == reqIndex ? way1Dirty_67 : _GEN_975; // @[DCache.scala 136:{22,22}]
  wire  _GEN_977 = 7'h44 == reqIndex ? way1Dirty_68 : _GEN_976; // @[DCache.scala 136:{22,22}]
  wire  _GEN_978 = 7'h45 == reqIndex ? way1Dirty_69 : _GEN_977; // @[DCache.scala 136:{22,22}]
  wire  _GEN_979 = 7'h46 == reqIndex ? way1Dirty_70 : _GEN_978; // @[DCache.scala 136:{22,22}]
  wire  _GEN_980 = 7'h47 == reqIndex ? way1Dirty_71 : _GEN_979; // @[DCache.scala 136:{22,22}]
  wire  _GEN_981 = 7'h48 == reqIndex ? way1Dirty_72 : _GEN_980; // @[DCache.scala 136:{22,22}]
  wire  _GEN_982 = 7'h49 == reqIndex ? way1Dirty_73 : _GEN_981; // @[DCache.scala 136:{22,22}]
  wire  _GEN_983 = 7'h4a == reqIndex ? way1Dirty_74 : _GEN_982; // @[DCache.scala 136:{22,22}]
  wire  _GEN_984 = 7'h4b == reqIndex ? way1Dirty_75 : _GEN_983; // @[DCache.scala 136:{22,22}]
  wire  _GEN_985 = 7'h4c == reqIndex ? way1Dirty_76 : _GEN_984; // @[DCache.scala 136:{22,22}]
  wire  _GEN_986 = 7'h4d == reqIndex ? way1Dirty_77 : _GEN_985; // @[DCache.scala 136:{22,22}]
  wire  _GEN_987 = 7'h4e == reqIndex ? way1Dirty_78 : _GEN_986; // @[DCache.scala 136:{22,22}]
  wire  _GEN_988 = 7'h4f == reqIndex ? way1Dirty_79 : _GEN_987; // @[DCache.scala 136:{22,22}]
  wire  _GEN_989 = 7'h50 == reqIndex ? way1Dirty_80 : _GEN_988; // @[DCache.scala 136:{22,22}]
  wire  _GEN_990 = 7'h51 == reqIndex ? way1Dirty_81 : _GEN_989; // @[DCache.scala 136:{22,22}]
  wire  _GEN_991 = 7'h52 == reqIndex ? way1Dirty_82 : _GEN_990; // @[DCache.scala 136:{22,22}]
  wire  _GEN_992 = 7'h53 == reqIndex ? way1Dirty_83 : _GEN_991; // @[DCache.scala 136:{22,22}]
  wire  _GEN_993 = 7'h54 == reqIndex ? way1Dirty_84 : _GEN_992; // @[DCache.scala 136:{22,22}]
  wire  _GEN_994 = 7'h55 == reqIndex ? way1Dirty_85 : _GEN_993; // @[DCache.scala 136:{22,22}]
  wire  _GEN_995 = 7'h56 == reqIndex ? way1Dirty_86 : _GEN_994; // @[DCache.scala 136:{22,22}]
  wire  _GEN_996 = 7'h57 == reqIndex ? way1Dirty_87 : _GEN_995; // @[DCache.scala 136:{22,22}]
  wire  _GEN_997 = 7'h58 == reqIndex ? way1Dirty_88 : _GEN_996; // @[DCache.scala 136:{22,22}]
  wire  _GEN_998 = 7'h59 == reqIndex ? way1Dirty_89 : _GEN_997; // @[DCache.scala 136:{22,22}]
  wire  _GEN_999 = 7'h5a == reqIndex ? way1Dirty_90 : _GEN_998; // @[DCache.scala 136:{22,22}]
  wire  _GEN_1000 = 7'h5b == reqIndex ? way1Dirty_91 : _GEN_999; // @[DCache.scala 136:{22,22}]
  wire  _GEN_1001 = 7'h5c == reqIndex ? way1Dirty_92 : _GEN_1000; // @[DCache.scala 136:{22,22}]
  wire  _GEN_1002 = 7'h5d == reqIndex ? way1Dirty_93 : _GEN_1001; // @[DCache.scala 136:{22,22}]
  wire  _GEN_1003 = 7'h5e == reqIndex ? way1Dirty_94 : _GEN_1002; // @[DCache.scala 136:{22,22}]
  wire  _GEN_1004 = 7'h5f == reqIndex ? way1Dirty_95 : _GEN_1003; // @[DCache.scala 136:{22,22}]
  wire  _GEN_1005 = 7'h60 == reqIndex ? way1Dirty_96 : _GEN_1004; // @[DCache.scala 136:{22,22}]
  wire  _GEN_1006 = 7'h61 == reqIndex ? way1Dirty_97 : _GEN_1005; // @[DCache.scala 136:{22,22}]
  wire  _GEN_1007 = 7'h62 == reqIndex ? way1Dirty_98 : _GEN_1006; // @[DCache.scala 136:{22,22}]
  wire  _GEN_1008 = 7'h63 == reqIndex ? way1Dirty_99 : _GEN_1007; // @[DCache.scala 136:{22,22}]
  wire  _GEN_1009 = 7'h64 == reqIndex ? way1Dirty_100 : _GEN_1008; // @[DCache.scala 136:{22,22}]
  wire  _GEN_1010 = 7'h65 == reqIndex ? way1Dirty_101 : _GEN_1009; // @[DCache.scala 136:{22,22}]
  wire  _GEN_1011 = 7'h66 == reqIndex ? way1Dirty_102 : _GEN_1010; // @[DCache.scala 136:{22,22}]
  wire  _GEN_1012 = 7'h67 == reqIndex ? way1Dirty_103 : _GEN_1011; // @[DCache.scala 136:{22,22}]
  wire  _GEN_1013 = 7'h68 == reqIndex ? way1Dirty_104 : _GEN_1012; // @[DCache.scala 136:{22,22}]
  wire  _GEN_1014 = 7'h69 == reqIndex ? way1Dirty_105 : _GEN_1013; // @[DCache.scala 136:{22,22}]
  wire  _GEN_1015 = 7'h6a == reqIndex ? way1Dirty_106 : _GEN_1014; // @[DCache.scala 136:{22,22}]
  wire  _GEN_1016 = 7'h6b == reqIndex ? way1Dirty_107 : _GEN_1015; // @[DCache.scala 136:{22,22}]
  wire  _GEN_1017 = 7'h6c == reqIndex ? way1Dirty_108 : _GEN_1016; // @[DCache.scala 136:{22,22}]
  wire  _GEN_1018 = 7'h6d == reqIndex ? way1Dirty_109 : _GEN_1017; // @[DCache.scala 136:{22,22}]
  wire  _GEN_1019 = 7'h6e == reqIndex ? way1Dirty_110 : _GEN_1018; // @[DCache.scala 136:{22,22}]
  wire  _GEN_1020 = 7'h6f == reqIndex ? way1Dirty_111 : _GEN_1019; // @[DCache.scala 136:{22,22}]
  wire  _GEN_1021 = 7'h70 == reqIndex ? way1Dirty_112 : _GEN_1020; // @[DCache.scala 136:{22,22}]
  wire  _GEN_1022 = 7'h71 == reqIndex ? way1Dirty_113 : _GEN_1021; // @[DCache.scala 136:{22,22}]
  wire  _GEN_1023 = 7'h72 == reqIndex ? way1Dirty_114 : _GEN_1022; // @[DCache.scala 136:{22,22}]
  wire  _GEN_1024 = 7'h73 == reqIndex ? way1Dirty_115 : _GEN_1023; // @[DCache.scala 136:{22,22}]
  wire  _GEN_1025 = 7'h74 == reqIndex ? way1Dirty_116 : _GEN_1024; // @[DCache.scala 136:{22,22}]
  wire  _GEN_1026 = 7'h75 == reqIndex ? way1Dirty_117 : _GEN_1025; // @[DCache.scala 136:{22,22}]
  wire  _GEN_1027 = 7'h76 == reqIndex ? way1Dirty_118 : _GEN_1026; // @[DCache.scala 136:{22,22}]
  wire  _GEN_1028 = 7'h77 == reqIndex ? way1Dirty_119 : _GEN_1027; // @[DCache.scala 136:{22,22}]
  wire  _GEN_1029 = 7'h78 == reqIndex ? way1Dirty_120 : _GEN_1028; // @[DCache.scala 136:{22,22}]
  wire  _GEN_1030 = 7'h79 == reqIndex ? way1Dirty_121 : _GEN_1029; // @[DCache.scala 136:{22,22}]
  wire  _GEN_1031 = 7'h7a == reqIndex ? way1Dirty_122 : _GEN_1030; // @[DCache.scala 136:{22,22}]
  wire  _GEN_1032 = 7'h7b == reqIndex ? way1Dirty_123 : _GEN_1031; // @[DCache.scala 136:{22,22}]
  wire  _GEN_1033 = 7'h7c == reqIndex ? way1Dirty_124 : _GEN_1032; // @[DCache.scala 136:{22,22}]
  wire  _GEN_1034 = 7'h7d == reqIndex ? way1Dirty_125 : _GEN_1033; // @[DCache.scala 136:{22,22}]
  wire  _GEN_1035 = 7'h7e == reqIndex ? way1Dirty_126 : _GEN_1034; // @[DCache.scala 136:{22,22}]
  wire  _GEN_1036 = 7'h7f == reqIndex ? way1Dirty_127 : _GEN_1035; // @[DCache.scala 136:{22,22}]
  wire  cacheDirtyEn = ~cacheLineWay ? _GEN_908 : _GEN_1036; // @[DCache.scala 136:22]
  wire [2:0] _GEN_3 = cacheDirtyEn ? 3'h3 : 3'h4; // @[DCache.scala 95:28 96:15 98:15]
  wire [2:0] _GEN_4 = io_out_data_ready ? 3'h4 : state; // @[DCache.scala 102:30 103:15 46:22]
  wire [2:0] _GEN_5 = io_out_data_ready ? 3'h5 : state; // @[DCache.scala 107:29 108:15 46:22]
  wire [2:0] _GEN_6 = 3'h6 == state ? 3'h0 : state; // @[DCache.scala 115:13 77:17 46:22]
  wire [2:0] _GEN_7 = 3'h5 == state ? 3'h6 : _GEN_6; // @[DCache.scala 112:15 77:17]
  wire [2:0] _GEN_8 = 3'h4 == state ? _GEN_5 : _GEN_7; // @[DCache.scala 77:17]
  wire [2:0] _GEN_9 = 3'h3 == state ? _GEN_4 : _GEN_8; // @[DCache.scala 77:17]
  wire  sHitEn = state == 3'h1; // @[DCache.scala 123:22]
  wire  _GEN_654 = 7'h1 == reqIndex ? way1Age_1 : way1Age_0; // @[DCache.scala 130:{53,53}]
  wire  _GEN_655 = 7'h2 == reqIndex ? way1Age_2 : _GEN_654; // @[DCache.scala 130:{53,53}]
  wire  _GEN_656 = 7'h3 == reqIndex ? way1Age_3 : _GEN_655; // @[DCache.scala 130:{53,53}]
  wire  _GEN_657 = 7'h4 == reqIndex ? way1Age_4 : _GEN_656; // @[DCache.scala 130:{53,53}]
  wire  _GEN_658 = 7'h5 == reqIndex ? way1Age_5 : _GEN_657; // @[DCache.scala 130:{53,53}]
  wire  _GEN_659 = 7'h6 == reqIndex ? way1Age_6 : _GEN_658; // @[DCache.scala 130:{53,53}]
  wire  _GEN_660 = 7'h7 == reqIndex ? way1Age_7 : _GEN_659; // @[DCache.scala 130:{53,53}]
  wire  _GEN_661 = 7'h8 == reqIndex ? way1Age_8 : _GEN_660; // @[DCache.scala 130:{53,53}]
  wire  _GEN_662 = 7'h9 == reqIndex ? way1Age_9 : _GEN_661; // @[DCache.scala 130:{53,53}]
  wire  _GEN_663 = 7'ha == reqIndex ? way1Age_10 : _GEN_662; // @[DCache.scala 130:{53,53}]
  wire  _GEN_664 = 7'hb == reqIndex ? way1Age_11 : _GEN_663; // @[DCache.scala 130:{53,53}]
  wire  _GEN_665 = 7'hc == reqIndex ? way1Age_12 : _GEN_664; // @[DCache.scala 130:{53,53}]
  wire  _GEN_666 = 7'hd == reqIndex ? way1Age_13 : _GEN_665; // @[DCache.scala 130:{53,53}]
  wire  _GEN_667 = 7'he == reqIndex ? way1Age_14 : _GEN_666; // @[DCache.scala 130:{53,53}]
  wire  _GEN_668 = 7'hf == reqIndex ? way1Age_15 : _GEN_667; // @[DCache.scala 130:{53,53}]
  wire  _GEN_669 = 7'h10 == reqIndex ? way1Age_16 : _GEN_668; // @[DCache.scala 130:{53,53}]
  wire  _GEN_670 = 7'h11 == reqIndex ? way1Age_17 : _GEN_669; // @[DCache.scala 130:{53,53}]
  wire  _GEN_671 = 7'h12 == reqIndex ? way1Age_18 : _GEN_670; // @[DCache.scala 130:{53,53}]
  wire  _GEN_672 = 7'h13 == reqIndex ? way1Age_19 : _GEN_671; // @[DCache.scala 130:{53,53}]
  wire  _GEN_673 = 7'h14 == reqIndex ? way1Age_20 : _GEN_672; // @[DCache.scala 130:{53,53}]
  wire  _GEN_674 = 7'h15 == reqIndex ? way1Age_21 : _GEN_673; // @[DCache.scala 130:{53,53}]
  wire  _GEN_675 = 7'h16 == reqIndex ? way1Age_22 : _GEN_674; // @[DCache.scala 130:{53,53}]
  wire  _GEN_676 = 7'h17 == reqIndex ? way1Age_23 : _GEN_675; // @[DCache.scala 130:{53,53}]
  wire  _GEN_677 = 7'h18 == reqIndex ? way1Age_24 : _GEN_676; // @[DCache.scala 130:{53,53}]
  wire  _GEN_678 = 7'h19 == reqIndex ? way1Age_25 : _GEN_677; // @[DCache.scala 130:{53,53}]
  wire  _GEN_679 = 7'h1a == reqIndex ? way1Age_26 : _GEN_678; // @[DCache.scala 130:{53,53}]
  wire  _GEN_680 = 7'h1b == reqIndex ? way1Age_27 : _GEN_679; // @[DCache.scala 130:{53,53}]
  wire  _GEN_681 = 7'h1c == reqIndex ? way1Age_28 : _GEN_680; // @[DCache.scala 130:{53,53}]
  wire  _GEN_682 = 7'h1d == reqIndex ? way1Age_29 : _GEN_681; // @[DCache.scala 130:{53,53}]
  wire  _GEN_683 = 7'h1e == reqIndex ? way1Age_30 : _GEN_682; // @[DCache.scala 130:{53,53}]
  wire  _GEN_684 = 7'h1f == reqIndex ? way1Age_31 : _GEN_683; // @[DCache.scala 130:{53,53}]
  wire  _GEN_685 = 7'h20 == reqIndex ? way1Age_32 : _GEN_684; // @[DCache.scala 130:{53,53}]
  wire  _GEN_686 = 7'h21 == reqIndex ? way1Age_33 : _GEN_685; // @[DCache.scala 130:{53,53}]
  wire  _GEN_687 = 7'h22 == reqIndex ? way1Age_34 : _GEN_686; // @[DCache.scala 130:{53,53}]
  wire  _GEN_688 = 7'h23 == reqIndex ? way1Age_35 : _GEN_687; // @[DCache.scala 130:{53,53}]
  wire  _GEN_689 = 7'h24 == reqIndex ? way1Age_36 : _GEN_688; // @[DCache.scala 130:{53,53}]
  wire  _GEN_690 = 7'h25 == reqIndex ? way1Age_37 : _GEN_689; // @[DCache.scala 130:{53,53}]
  wire  _GEN_691 = 7'h26 == reqIndex ? way1Age_38 : _GEN_690; // @[DCache.scala 130:{53,53}]
  wire  _GEN_692 = 7'h27 == reqIndex ? way1Age_39 : _GEN_691; // @[DCache.scala 130:{53,53}]
  wire  _GEN_693 = 7'h28 == reqIndex ? way1Age_40 : _GEN_692; // @[DCache.scala 130:{53,53}]
  wire  _GEN_694 = 7'h29 == reqIndex ? way1Age_41 : _GEN_693; // @[DCache.scala 130:{53,53}]
  wire  _GEN_695 = 7'h2a == reqIndex ? way1Age_42 : _GEN_694; // @[DCache.scala 130:{53,53}]
  wire  _GEN_696 = 7'h2b == reqIndex ? way1Age_43 : _GEN_695; // @[DCache.scala 130:{53,53}]
  wire  _GEN_697 = 7'h2c == reqIndex ? way1Age_44 : _GEN_696; // @[DCache.scala 130:{53,53}]
  wire  _GEN_698 = 7'h2d == reqIndex ? way1Age_45 : _GEN_697; // @[DCache.scala 130:{53,53}]
  wire  _GEN_699 = 7'h2e == reqIndex ? way1Age_46 : _GEN_698; // @[DCache.scala 130:{53,53}]
  wire  _GEN_700 = 7'h2f == reqIndex ? way1Age_47 : _GEN_699; // @[DCache.scala 130:{53,53}]
  wire  _GEN_701 = 7'h30 == reqIndex ? way1Age_48 : _GEN_700; // @[DCache.scala 130:{53,53}]
  wire  _GEN_702 = 7'h31 == reqIndex ? way1Age_49 : _GEN_701; // @[DCache.scala 130:{53,53}]
  wire  _GEN_703 = 7'h32 == reqIndex ? way1Age_50 : _GEN_702; // @[DCache.scala 130:{53,53}]
  wire  _GEN_704 = 7'h33 == reqIndex ? way1Age_51 : _GEN_703; // @[DCache.scala 130:{53,53}]
  wire  _GEN_705 = 7'h34 == reqIndex ? way1Age_52 : _GEN_704; // @[DCache.scala 130:{53,53}]
  wire  _GEN_706 = 7'h35 == reqIndex ? way1Age_53 : _GEN_705; // @[DCache.scala 130:{53,53}]
  wire  _GEN_707 = 7'h36 == reqIndex ? way1Age_54 : _GEN_706; // @[DCache.scala 130:{53,53}]
  wire  _GEN_708 = 7'h37 == reqIndex ? way1Age_55 : _GEN_707; // @[DCache.scala 130:{53,53}]
  wire  _GEN_709 = 7'h38 == reqIndex ? way1Age_56 : _GEN_708; // @[DCache.scala 130:{53,53}]
  wire  _GEN_710 = 7'h39 == reqIndex ? way1Age_57 : _GEN_709; // @[DCache.scala 130:{53,53}]
  wire  _GEN_711 = 7'h3a == reqIndex ? way1Age_58 : _GEN_710; // @[DCache.scala 130:{53,53}]
  wire  _GEN_712 = 7'h3b == reqIndex ? way1Age_59 : _GEN_711; // @[DCache.scala 130:{53,53}]
  wire  _GEN_713 = 7'h3c == reqIndex ? way1Age_60 : _GEN_712; // @[DCache.scala 130:{53,53}]
  wire  _GEN_714 = 7'h3d == reqIndex ? way1Age_61 : _GEN_713; // @[DCache.scala 130:{53,53}]
  wire  _GEN_715 = 7'h3e == reqIndex ? way1Age_62 : _GEN_714; // @[DCache.scala 130:{53,53}]
  wire  _GEN_716 = 7'h3f == reqIndex ? way1Age_63 : _GEN_715; // @[DCache.scala 130:{53,53}]
  wire  _GEN_717 = 7'h40 == reqIndex ? way1Age_64 : _GEN_716; // @[DCache.scala 130:{53,53}]
  wire  _GEN_718 = 7'h41 == reqIndex ? way1Age_65 : _GEN_717; // @[DCache.scala 130:{53,53}]
  wire  _GEN_719 = 7'h42 == reqIndex ? way1Age_66 : _GEN_718; // @[DCache.scala 130:{53,53}]
  wire  _GEN_720 = 7'h43 == reqIndex ? way1Age_67 : _GEN_719; // @[DCache.scala 130:{53,53}]
  wire  _GEN_721 = 7'h44 == reqIndex ? way1Age_68 : _GEN_720; // @[DCache.scala 130:{53,53}]
  wire  _GEN_722 = 7'h45 == reqIndex ? way1Age_69 : _GEN_721; // @[DCache.scala 130:{53,53}]
  wire  _GEN_723 = 7'h46 == reqIndex ? way1Age_70 : _GEN_722; // @[DCache.scala 130:{53,53}]
  wire  _GEN_724 = 7'h47 == reqIndex ? way1Age_71 : _GEN_723; // @[DCache.scala 130:{53,53}]
  wire  _GEN_725 = 7'h48 == reqIndex ? way1Age_72 : _GEN_724; // @[DCache.scala 130:{53,53}]
  wire  _GEN_726 = 7'h49 == reqIndex ? way1Age_73 : _GEN_725; // @[DCache.scala 130:{53,53}]
  wire  _GEN_727 = 7'h4a == reqIndex ? way1Age_74 : _GEN_726; // @[DCache.scala 130:{53,53}]
  wire  _GEN_728 = 7'h4b == reqIndex ? way1Age_75 : _GEN_727; // @[DCache.scala 130:{53,53}]
  wire  _GEN_729 = 7'h4c == reqIndex ? way1Age_76 : _GEN_728; // @[DCache.scala 130:{53,53}]
  wire  _GEN_730 = 7'h4d == reqIndex ? way1Age_77 : _GEN_729; // @[DCache.scala 130:{53,53}]
  wire  _GEN_731 = 7'h4e == reqIndex ? way1Age_78 : _GEN_730; // @[DCache.scala 130:{53,53}]
  wire  _GEN_732 = 7'h4f == reqIndex ? way1Age_79 : _GEN_731; // @[DCache.scala 130:{53,53}]
  wire  _GEN_733 = 7'h50 == reqIndex ? way1Age_80 : _GEN_732; // @[DCache.scala 130:{53,53}]
  wire  _GEN_734 = 7'h51 == reqIndex ? way1Age_81 : _GEN_733; // @[DCache.scala 130:{53,53}]
  wire  _GEN_735 = 7'h52 == reqIndex ? way1Age_82 : _GEN_734; // @[DCache.scala 130:{53,53}]
  wire  _GEN_736 = 7'h53 == reqIndex ? way1Age_83 : _GEN_735; // @[DCache.scala 130:{53,53}]
  wire  _GEN_737 = 7'h54 == reqIndex ? way1Age_84 : _GEN_736; // @[DCache.scala 130:{53,53}]
  wire  _GEN_738 = 7'h55 == reqIndex ? way1Age_85 : _GEN_737; // @[DCache.scala 130:{53,53}]
  wire  _GEN_739 = 7'h56 == reqIndex ? way1Age_86 : _GEN_738; // @[DCache.scala 130:{53,53}]
  wire  _GEN_740 = 7'h57 == reqIndex ? way1Age_87 : _GEN_739; // @[DCache.scala 130:{53,53}]
  wire  _GEN_741 = 7'h58 == reqIndex ? way1Age_88 : _GEN_740; // @[DCache.scala 130:{53,53}]
  wire  _GEN_742 = 7'h59 == reqIndex ? way1Age_89 : _GEN_741; // @[DCache.scala 130:{53,53}]
  wire  _GEN_743 = 7'h5a == reqIndex ? way1Age_90 : _GEN_742; // @[DCache.scala 130:{53,53}]
  wire  _GEN_744 = 7'h5b == reqIndex ? way1Age_91 : _GEN_743; // @[DCache.scala 130:{53,53}]
  wire  _GEN_745 = 7'h5c == reqIndex ? way1Age_92 : _GEN_744; // @[DCache.scala 130:{53,53}]
  wire  _GEN_746 = 7'h5d == reqIndex ? way1Age_93 : _GEN_745; // @[DCache.scala 130:{53,53}]
  wire  _GEN_747 = 7'h5e == reqIndex ? way1Age_94 : _GEN_746; // @[DCache.scala 130:{53,53}]
  wire  _GEN_748 = 7'h5f == reqIndex ? way1Age_95 : _GEN_747; // @[DCache.scala 130:{53,53}]
  wire  _GEN_749 = 7'h60 == reqIndex ? way1Age_96 : _GEN_748; // @[DCache.scala 130:{53,53}]
  wire  _GEN_750 = 7'h61 == reqIndex ? way1Age_97 : _GEN_749; // @[DCache.scala 130:{53,53}]
  wire  _GEN_751 = 7'h62 == reqIndex ? way1Age_98 : _GEN_750; // @[DCache.scala 130:{53,53}]
  wire  _GEN_752 = 7'h63 == reqIndex ? way1Age_99 : _GEN_751; // @[DCache.scala 130:{53,53}]
  wire  _GEN_753 = 7'h64 == reqIndex ? way1Age_100 : _GEN_752; // @[DCache.scala 130:{53,53}]
  wire  _GEN_754 = 7'h65 == reqIndex ? way1Age_101 : _GEN_753; // @[DCache.scala 130:{53,53}]
  wire  _GEN_755 = 7'h66 == reqIndex ? way1Age_102 : _GEN_754; // @[DCache.scala 130:{53,53}]
  wire  _GEN_756 = 7'h67 == reqIndex ? way1Age_103 : _GEN_755; // @[DCache.scala 130:{53,53}]
  wire  _GEN_757 = 7'h68 == reqIndex ? way1Age_104 : _GEN_756; // @[DCache.scala 130:{53,53}]
  wire  _GEN_758 = 7'h69 == reqIndex ? way1Age_105 : _GEN_757; // @[DCache.scala 130:{53,53}]
  wire  _GEN_759 = 7'h6a == reqIndex ? way1Age_106 : _GEN_758; // @[DCache.scala 130:{53,53}]
  wire  _GEN_760 = 7'h6b == reqIndex ? way1Age_107 : _GEN_759; // @[DCache.scala 130:{53,53}]
  wire  _GEN_761 = 7'h6c == reqIndex ? way1Age_108 : _GEN_760; // @[DCache.scala 130:{53,53}]
  wire  _GEN_762 = 7'h6d == reqIndex ? way1Age_109 : _GEN_761; // @[DCache.scala 130:{53,53}]
  wire  _GEN_763 = 7'h6e == reqIndex ? way1Age_110 : _GEN_762; // @[DCache.scala 130:{53,53}]
  wire  _GEN_764 = 7'h6f == reqIndex ? way1Age_111 : _GEN_763; // @[DCache.scala 130:{53,53}]
  wire  _GEN_765 = 7'h70 == reqIndex ? way1Age_112 : _GEN_764; // @[DCache.scala 130:{53,53}]
  wire  _GEN_766 = 7'h71 == reqIndex ? way1Age_113 : _GEN_765; // @[DCache.scala 130:{53,53}]
  wire  _GEN_767 = 7'h72 == reqIndex ? way1Age_114 : _GEN_766; // @[DCache.scala 130:{53,53}]
  wire  _GEN_768 = 7'h73 == reqIndex ? way1Age_115 : _GEN_767; // @[DCache.scala 130:{53,53}]
  wire  _GEN_769 = 7'h74 == reqIndex ? way1Age_116 : _GEN_768; // @[DCache.scala 130:{53,53}]
  wire  _GEN_770 = 7'h75 == reqIndex ? way1Age_117 : _GEN_769; // @[DCache.scala 130:{53,53}]
  wire  _GEN_771 = 7'h76 == reqIndex ? way1Age_118 : _GEN_770; // @[DCache.scala 130:{53,53}]
  wire  _GEN_772 = 7'h77 == reqIndex ? way1Age_119 : _GEN_771; // @[DCache.scala 130:{53,53}]
  wire  _GEN_773 = 7'h78 == reqIndex ? way1Age_120 : _GEN_772; // @[DCache.scala 130:{53,53}]
  wire  _GEN_774 = 7'h79 == reqIndex ? way1Age_121 : _GEN_773; // @[DCache.scala 130:{53,53}]
  wire  _GEN_775 = 7'h7a == reqIndex ? way1Age_122 : _GEN_774; // @[DCache.scala 130:{53,53}]
  wire  _GEN_776 = 7'h7b == reqIndex ? way1Age_123 : _GEN_775; // @[DCache.scala 130:{53,53}]
  wire  _GEN_777 = 7'h7c == reqIndex ? way1Age_124 : _GEN_776; // @[DCache.scala 130:{53,53}]
  wire  _GEN_778 = 7'h7d == reqIndex ? way1Age_125 : _GEN_777; // @[DCache.scala 130:{53,53}]
  wire  _GEN_779 = 7'h7e == reqIndex ? way1Age_126 : _GEN_778; // @[DCache.scala 130:{53,53}]
  wire  _GEN_780 = 7'h7f == reqIndex ? way1Age_127 : _GEN_779; // @[DCache.scala 130:{53,53}]
  wire  ageWay1En = _ageWay0En_T & ~_GEN_780; // @[DCache.scala 130:31]
  wire [7:0] _cacheIndex_T_1 = {1'h0,reqIndex}; // @[Cat.scala 31:58]
  wire [7:0] _cacheIndex_T_2 = {1'h1,reqIndex}; // @[Cat.scala 31:58]
  wire  sWriteEn = state == 3'h3; // @[DCache.scala 138:24]
  wire  sReadEn = state == 3'h4; // @[DCache.scala 140:24]
  wire  sCacheWEn = state == 3'h5; // @[DCache.scala 142:26]
  wire [127:0] cacheRData = req_Q;
  wire [63:0] valid_data = reqOff[3] ? cacheRData[127:64] : cacheRData[63:0]; // @[DCache.scala 147:23]
  wire [63:0] inDataWT = reqOff[3] ? io_dmem_data_write[127:64] : io_dmem_data_write[63:0]; // @[DCache.scala 148:23]
  wire [63:0] _cacheWDataT_T_3 = {valid_data[63:8],inDataWT[7:0]}; // @[Cat.scala 31:58]
  wire [63:0] _cacheWDataT_T_7 = {valid_data[63:16],inDataWT[15:8],valid_data[7:0]}; // @[Cat.scala 31:58]
  wire [63:0] _cacheWDataT_T_11 = {valid_data[63:24],inDataWT[23:16],valid_data[15:0]}; // @[Cat.scala 31:58]
  wire [63:0] _cacheWDataT_T_15 = {valid_data[63:32],inDataWT[31:24],valid_data[23:0]}; // @[Cat.scala 31:58]
  wire [63:0] _cacheWDataT_T_19 = {valid_data[63:40],inDataWT[39:32],valid_data[31:0]}; // @[Cat.scala 31:58]
  wire [63:0] _cacheWDataT_T_23 = {valid_data[63:48],inDataWT[47:40],valid_data[39:0]}; // @[Cat.scala 31:58]
  wire [63:0] _cacheWDataT_T_27 = {valid_data[63:56],inDataWT[55:48],valid_data[47:0]}; // @[Cat.scala 31:58]
  wire [63:0] _cacheWDataT_T_30 = {inDataWT[63:56],valid_data[55:0]}; // @[Cat.scala 31:58]
  wire [63:0] _cacheWDataT_T_32 = 3'h1 == reqOff[2:0] ? _cacheWDataT_T_7 : _cacheWDataT_T_3; // @[Mux.scala 81:58]
  wire [63:0] _cacheWDataT_T_34 = 3'h2 == reqOff[2:0] ? _cacheWDataT_T_11 : _cacheWDataT_T_32; // @[Mux.scala 81:58]
  wire [63:0] _cacheWDataT_T_36 = 3'h3 == reqOff[2:0] ? _cacheWDataT_T_15 : _cacheWDataT_T_34; // @[Mux.scala 81:58]
  wire [63:0] _cacheWDataT_T_38 = 3'h4 == reqOff[2:0] ? _cacheWDataT_T_19 : _cacheWDataT_T_36; // @[Mux.scala 81:58]
  wire [63:0] _cacheWDataT_T_40 = 3'h5 == reqOff[2:0] ? _cacheWDataT_T_23 : _cacheWDataT_T_38; // @[Mux.scala 81:58]
  wire [63:0] _cacheWDataT_T_42 = 3'h6 == reqOff[2:0] ? _cacheWDataT_T_27 : _cacheWDataT_T_40; // @[Mux.scala 81:58]
  wire [63:0] _cacheWDataT_T_44 = 3'h7 == reqOff[2:0] ? _cacheWDataT_T_30 : _cacheWDataT_T_42; // @[Mux.scala 81:58]
  wire [63:0] _cacheWDataT_T_48 = {valid_data[63:16],inDataWT[15:0]}; // @[Cat.scala 31:58]
  wire [63:0] _cacheWDataT_T_52 = {valid_data[63:32],inDataWT[31:16],valid_data[15:0]}; // @[Cat.scala 31:58]
  wire [63:0] _cacheWDataT_T_56 = {valid_data[63:48],inDataWT[47:32],valid_data[31:0]}; // @[Cat.scala 31:58]
  wire [63:0] _cacheWDataT_T_59 = {inDataWT[63:48],valid_data[47:0]}; // @[Cat.scala 31:58]
  wire [63:0] _cacheWDataT_T_61 = 2'h1 == reqOff[2:1] ? _cacheWDataT_T_52 : _cacheWDataT_T_48; // @[Mux.scala 81:58]
  wire [63:0] _cacheWDataT_T_63 = 2'h2 == reqOff[2:1] ? _cacheWDataT_T_56 : _cacheWDataT_T_61; // @[Mux.scala 81:58]
  wire [63:0] _cacheWDataT_T_65 = 2'h3 == reqOff[2:1] ? _cacheWDataT_T_59 : _cacheWDataT_T_63; // @[Mux.scala 81:58]
  wire [63:0] _cacheWDataT_T_69 = {valid_data[63:32],inDataWT[31:0]}; // @[Cat.scala 31:58]
  wire [63:0] _cacheWDataT_T_72 = {inDataWT[63:32],valid_data[31:0]}; // @[Cat.scala 31:58]
  wire [63:0] _cacheWDataT_T_74 = reqOff[2] ? _cacheWDataT_T_72 : _cacheWDataT_T_69; // @[Mux.scala 81:58]
  wire [63:0] _cacheWDataT_T_76 = 2'h1 == io_dmem_data_size ? _cacheWDataT_T_65 : _cacheWDataT_T_44; // @[Mux.scala 81:58]
  wire [63:0] _cacheWDataT_T_78 = 2'h2 == io_dmem_data_size ? _cacheWDataT_T_74 : _cacheWDataT_T_76; // @[Mux.scala 81:58]
  wire [63:0] cacheWDataT = 2'h3 == io_dmem_data_size ? inDataWT : _cacheWDataT_T_78; // @[Mux.scala 81:58]
  wire [127:0] _cacheWData_T_1 = {cacheWDataT,64'h0}; // @[Cat.scala 31:58]
  wire [127:0] _cacheWData_T_2 = {64'h0,cacheWDataT}; // @[Cat.scala 31:58]
  wire [127:0] cacheWData = reqOff[3] ? _cacheWData_T_1 : _cacheWData_T_2; // @[DCache.scala 172:23]
  wire  _valid_WEn_T = sReadEn & io_out_data_ready; // @[DCache.scala 175:40]
  wire [127:0] _valid_WData_T_1 = io_dmem_data_req ? cacheWData : io_out_data_read; // @[DCache.scala 177:22]
  wire [127:0] _valid_BWEn_T_1 = io_dmem_data_req ? valid_strb : 128'hffffffffffffffffffffffffffffffff; // @[DCache.scala 179:22]
  wire  _T_9 = sCacheWEn & io_dmem_data_req; // @[DCache.scala 183:20]
  wire  _GEN_4749 = 7'h0 == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1037 = 7'h0 == reqIndex | way0Dirty_0; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4750 = 7'h1 == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1038 = 7'h1 == reqIndex | way0Dirty_1; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4751 = 7'h2 == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1039 = 7'h2 == reqIndex | way0Dirty_2; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4752 = 7'h3 == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1040 = 7'h3 == reqIndex | way0Dirty_3; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4753 = 7'h4 == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1041 = 7'h4 == reqIndex | way0Dirty_4; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4754 = 7'h5 == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1042 = 7'h5 == reqIndex | way0Dirty_5; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4755 = 7'h6 == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1043 = 7'h6 == reqIndex | way0Dirty_6; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4756 = 7'h7 == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1044 = 7'h7 == reqIndex | way0Dirty_7; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4757 = 7'h8 == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1045 = 7'h8 == reqIndex | way0Dirty_8; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4758 = 7'h9 == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1046 = 7'h9 == reqIndex | way0Dirty_9; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4759 = 7'ha == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1047 = 7'ha == reqIndex | way0Dirty_10; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4760 = 7'hb == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1048 = 7'hb == reqIndex | way0Dirty_11; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4761 = 7'hc == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1049 = 7'hc == reqIndex | way0Dirty_12; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4762 = 7'hd == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1050 = 7'hd == reqIndex | way0Dirty_13; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4763 = 7'he == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1051 = 7'he == reqIndex | way0Dirty_14; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4764 = 7'hf == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1052 = 7'hf == reqIndex | way0Dirty_15; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4765 = 7'h10 == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1053 = 7'h10 == reqIndex | way0Dirty_16; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4766 = 7'h11 == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1054 = 7'h11 == reqIndex | way0Dirty_17; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4767 = 7'h12 == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1055 = 7'h12 == reqIndex | way0Dirty_18; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4768 = 7'h13 == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1056 = 7'h13 == reqIndex | way0Dirty_19; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4769 = 7'h14 == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1057 = 7'h14 == reqIndex | way0Dirty_20; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4770 = 7'h15 == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1058 = 7'h15 == reqIndex | way0Dirty_21; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4771 = 7'h16 == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1059 = 7'h16 == reqIndex | way0Dirty_22; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4772 = 7'h17 == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1060 = 7'h17 == reqIndex | way0Dirty_23; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4773 = 7'h18 == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1061 = 7'h18 == reqIndex | way0Dirty_24; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4774 = 7'h19 == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1062 = 7'h19 == reqIndex | way0Dirty_25; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4775 = 7'h1a == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1063 = 7'h1a == reqIndex | way0Dirty_26; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4776 = 7'h1b == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1064 = 7'h1b == reqIndex | way0Dirty_27; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4777 = 7'h1c == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1065 = 7'h1c == reqIndex | way0Dirty_28; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4778 = 7'h1d == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1066 = 7'h1d == reqIndex | way0Dirty_29; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4779 = 7'h1e == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1067 = 7'h1e == reqIndex | way0Dirty_30; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4780 = 7'h1f == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1068 = 7'h1f == reqIndex | way0Dirty_31; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4781 = 7'h20 == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1069 = 7'h20 == reqIndex | way0Dirty_32; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4782 = 7'h21 == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1070 = 7'h21 == reqIndex | way0Dirty_33; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4783 = 7'h22 == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1071 = 7'h22 == reqIndex | way0Dirty_34; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4784 = 7'h23 == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1072 = 7'h23 == reqIndex | way0Dirty_35; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4785 = 7'h24 == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1073 = 7'h24 == reqIndex | way0Dirty_36; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4786 = 7'h25 == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1074 = 7'h25 == reqIndex | way0Dirty_37; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4787 = 7'h26 == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1075 = 7'h26 == reqIndex | way0Dirty_38; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4788 = 7'h27 == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1076 = 7'h27 == reqIndex | way0Dirty_39; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4789 = 7'h28 == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1077 = 7'h28 == reqIndex | way0Dirty_40; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4790 = 7'h29 == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1078 = 7'h29 == reqIndex | way0Dirty_41; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4791 = 7'h2a == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1079 = 7'h2a == reqIndex | way0Dirty_42; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4792 = 7'h2b == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1080 = 7'h2b == reqIndex | way0Dirty_43; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4793 = 7'h2c == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1081 = 7'h2c == reqIndex | way0Dirty_44; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4794 = 7'h2d == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1082 = 7'h2d == reqIndex | way0Dirty_45; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4795 = 7'h2e == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1083 = 7'h2e == reqIndex | way0Dirty_46; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4796 = 7'h2f == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1084 = 7'h2f == reqIndex | way0Dirty_47; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4797 = 7'h30 == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1085 = 7'h30 == reqIndex | way0Dirty_48; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4798 = 7'h31 == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1086 = 7'h31 == reqIndex | way0Dirty_49; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4799 = 7'h32 == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1087 = 7'h32 == reqIndex | way0Dirty_50; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4800 = 7'h33 == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1088 = 7'h33 == reqIndex | way0Dirty_51; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4801 = 7'h34 == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1089 = 7'h34 == reqIndex | way0Dirty_52; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4802 = 7'h35 == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1090 = 7'h35 == reqIndex | way0Dirty_53; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4803 = 7'h36 == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1091 = 7'h36 == reqIndex | way0Dirty_54; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4804 = 7'h37 == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1092 = 7'h37 == reqIndex | way0Dirty_55; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4805 = 7'h38 == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1093 = 7'h38 == reqIndex | way0Dirty_56; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4806 = 7'h39 == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1094 = 7'h39 == reqIndex | way0Dirty_57; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4807 = 7'h3a == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1095 = 7'h3a == reqIndex | way0Dirty_58; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4808 = 7'h3b == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1096 = 7'h3b == reqIndex | way0Dirty_59; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4809 = 7'h3c == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1097 = 7'h3c == reqIndex | way0Dirty_60; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4810 = 7'h3d == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1098 = 7'h3d == reqIndex | way0Dirty_61; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4811 = 7'h3e == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1099 = 7'h3e == reqIndex | way0Dirty_62; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4812 = 7'h3f == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1100 = 7'h3f == reqIndex | way0Dirty_63; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4813 = 7'h40 == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1101 = 7'h40 == reqIndex | way0Dirty_64; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4814 = 7'h41 == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1102 = 7'h41 == reqIndex | way0Dirty_65; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4815 = 7'h42 == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1103 = 7'h42 == reqIndex | way0Dirty_66; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4816 = 7'h43 == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1104 = 7'h43 == reqIndex | way0Dirty_67; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4817 = 7'h44 == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1105 = 7'h44 == reqIndex | way0Dirty_68; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4818 = 7'h45 == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1106 = 7'h45 == reqIndex | way0Dirty_69; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4819 = 7'h46 == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1107 = 7'h46 == reqIndex | way0Dirty_70; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4820 = 7'h47 == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1108 = 7'h47 == reqIndex | way0Dirty_71; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4821 = 7'h48 == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1109 = 7'h48 == reqIndex | way0Dirty_72; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4822 = 7'h49 == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1110 = 7'h49 == reqIndex | way0Dirty_73; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4823 = 7'h4a == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1111 = 7'h4a == reqIndex | way0Dirty_74; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4824 = 7'h4b == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1112 = 7'h4b == reqIndex | way0Dirty_75; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4825 = 7'h4c == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1113 = 7'h4c == reqIndex | way0Dirty_76; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4826 = 7'h4d == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1114 = 7'h4d == reqIndex | way0Dirty_77; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4827 = 7'h4e == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1115 = 7'h4e == reqIndex | way0Dirty_78; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4828 = 7'h4f == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1116 = 7'h4f == reqIndex | way0Dirty_79; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4829 = 7'h50 == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1117 = 7'h50 == reqIndex | way0Dirty_80; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4830 = 7'h51 == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1118 = 7'h51 == reqIndex | way0Dirty_81; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4831 = 7'h52 == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1119 = 7'h52 == reqIndex | way0Dirty_82; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4832 = 7'h53 == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1120 = 7'h53 == reqIndex | way0Dirty_83; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4833 = 7'h54 == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1121 = 7'h54 == reqIndex | way0Dirty_84; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4834 = 7'h55 == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1122 = 7'h55 == reqIndex | way0Dirty_85; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4835 = 7'h56 == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1123 = 7'h56 == reqIndex | way0Dirty_86; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4836 = 7'h57 == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1124 = 7'h57 == reqIndex | way0Dirty_87; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4837 = 7'h58 == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1125 = 7'h58 == reqIndex | way0Dirty_88; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4838 = 7'h59 == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1126 = 7'h59 == reqIndex | way0Dirty_89; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4839 = 7'h5a == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1127 = 7'h5a == reqIndex | way0Dirty_90; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4840 = 7'h5b == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1128 = 7'h5b == reqIndex | way0Dirty_91; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4841 = 7'h5c == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1129 = 7'h5c == reqIndex | way0Dirty_92; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4842 = 7'h5d == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1130 = 7'h5d == reqIndex | way0Dirty_93; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4843 = 7'h5e == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1131 = 7'h5e == reqIndex | way0Dirty_94; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4844 = 7'h5f == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1132 = 7'h5f == reqIndex | way0Dirty_95; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4845 = 7'h60 == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1133 = 7'h60 == reqIndex | way0Dirty_96; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4846 = 7'h61 == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1134 = 7'h61 == reqIndex | way0Dirty_97; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4847 = 7'h62 == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1135 = 7'h62 == reqIndex | way0Dirty_98; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4848 = 7'h63 == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1136 = 7'h63 == reqIndex | way0Dirty_99; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4849 = 7'h64 == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1137 = 7'h64 == reqIndex | way0Dirty_100; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4850 = 7'h65 == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1138 = 7'h65 == reqIndex | way0Dirty_101; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4851 = 7'h66 == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1139 = 7'h66 == reqIndex | way0Dirty_102; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4852 = 7'h67 == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1140 = 7'h67 == reqIndex | way0Dirty_103; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4853 = 7'h68 == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1141 = 7'h68 == reqIndex | way0Dirty_104; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4854 = 7'h69 == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1142 = 7'h69 == reqIndex | way0Dirty_105; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4855 = 7'h6a == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1143 = 7'h6a == reqIndex | way0Dirty_106; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4856 = 7'h6b == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1144 = 7'h6b == reqIndex | way0Dirty_107; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4857 = 7'h6c == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1145 = 7'h6c == reqIndex | way0Dirty_108; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4858 = 7'h6d == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1146 = 7'h6d == reqIndex | way0Dirty_109; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4859 = 7'h6e == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1147 = 7'h6e == reqIndex | way0Dirty_110; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4860 = 7'h6f == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1148 = 7'h6f == reqIndex | way0Dirty_111; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4861 = 7'h70 == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1149 = 7'h70 == reqIndex | way0Dirty_112; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4862 = 7'h71 == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1150 = 7'h71 == reqIndex | way0Dirty_113; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4863 = 7'h72 == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1151 = 7'h72 == reqIndex | way0Dirty_114; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4864 = 7'h73 == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1152 = 7'h73 == reqIndex | way0Dirty_115; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4865 = 7'h74 == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1153 = 7'h74 == reqIndex | way0Dirty_116; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4866 = 7'h75 == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1154 = 7'h75 == reqIndex | way0Dirty_117; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4867 = 7'h76 == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1155 = 7'h76 == reqIndex | way0Dirty_118; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4868 = 7'h77 == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1156 = 7'h77 == reqIndex | way0Dirty_119; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4869 = 7'h78 == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1157 = 7'h78 == reqIndex | way0Dirty_120; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4870 = 7'h79 == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1158 = 7'h79 == reqIndex | way0Dirty_121; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4871 = 7'h7a == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1159 = 7'h7a == reqIndex | way0Dirty_122; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4872 = 7'h7b == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1160 = 7'h7b == reqIndex | way0Dirty_123; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4873 = 7'h7c == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1161 = 7'h7c == reqIndex | way0Dirty_124; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4874 = 7'h7d == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1162 = 7'h7d == reqIndex | way0Dirty_125; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4875 = 7'h7e == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1163 = 7'h7e == reqIndex | way0Dirty_126; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_4876 = 7'h7f == reqIndex; // @[DCache.scala 184:{27,27} 37:26]
  wire  _GEN_1164 = 7'h7f == reqIndex | way0Dirty_127; // @[DCache.scala 184:{27,27} 37:26]
  wire  _T_10 = sWriteEn & io_out_data_ready; // @[DCache.scala 185:26]
  wire  _GEN_1165 = 7'h0 == reqIndex ? 1'h0 : way0Dirty_0; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1166 = 7'h1 == reqIndex ? 1'h0 : way0Dirty_1; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1167 = 7'h2 == reqIndex ? 1'h0 : way0Dirty_2; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1168 = 7'h3 == reqIndex ? 1'h0 : way0Dirty_3; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1169 = 7'h4 == reqIndex ? 1'h0 : way0Dirty_4; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1170 = 7'h5 == reqIndex ? 1'h0 : way0Dirty_5; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1171 = 7'h6 == reqIndex ? 1'h0 : way0Dirty_6; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1172 = 7'h7 == reqIndex ? 1'h0 : way0Dirty_7; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1173 = 7'h8 == reqIndex ? 1'h0 : way0Dirty_8; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1174 = 7'h9 == reqIndex ? 1'h0 : way0Dirty_9; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1175 = 7'ha == reqIndex ? 1'h0 : way0Dirty_10; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1176 = 7'hb == reqIndex ? 1'h0 : way0Dirty_11; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1177 = 7'hc == reqIndex ? 1'h0 : way0Dirty_12; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1178 = 7'hd == reqIndex ? 1'h0 : way0Dirty_13; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1179 = 7'he == reqIndex ? 1'h0 : way0Dirty_14; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1180 = 7'hf == reqIndex ? 1'h0 : way0Dirty_15; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1181 = 7'h10 == reqIndex ? 1'h0 : way0Dirty_16; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1182 = 7'h11 == reqIndex ? 1'h0 : way0Dirty_17; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1183 = 7'h12 == reqIndex ? 1'h0 : way0Dirty_18; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1184 = 7'h13 == reqIndex ? 1'h0 : way0Dirty_19; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1185 = 7'h14 == reqIndex ? 1'h0 : way0Dirty_20; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1186 = 7'h15 == reqIndex ? 1'h0 : way0Dirty_21; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1187 = 7'h16 == reqIndex ? 1'h0 : way0Dirty_22; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1188 = 7'h17 == reqIndex ? 1'h0 : way0Dirty_23; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1189 = 7'h18 == reqIndex ? 1'h0 : way0Dirty_24; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1190 = 7'h19 == reqIndex ? 1'h0 : way0Dirty_25; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1191 = 7'h1a == reqIndex ? 1'h0 : way0Dirty_26; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1192 = 7'h1b == reqIndex ? 1'h0 : way0Dirty_27; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1193 = 7'h1c == reqIndex ? 1'h0 : way0Dirty_28; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1194 = 7'h1d == reqIndex ? 1'h0 : way0Dirty_29; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1195 = 7'h1e == reqIndex ? 1'h0 : way0Dirty_30; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1196 = 7'h1f == reqIndex ? 1'h0 : way0Dirty_31; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1197 = 7'h20 == reqIndex ? 1'h0 : way0Dirty_32; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1198 = 7'h21 == reqIndex ? 1'h0 : way0Dirty_33; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1199 = 7'h22 == reqIndex ? 1'h0 : way0Dirty_34; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1200 = 7'h23 == reqIndex ? 1'h0 : way0Dirty_35; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1201 = 7'h24 == reqIndex ? 1'h0 : way0Dirty_36; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1202 = 7'h25 == reqIndex ? 1'h0 : way0Dirty_37; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1203 = 7'h26 == reqIndex ? 1'h0 : way0Dirty_38; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1204 = 7'h27 == reqIndex ? 1'h0 : way0Dirty_39; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1205 = 7'h28 == reqIndex ? 1'h0 : way0Dirty_40; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1206 = 7'h29 == reqIndex ? 1'h0 : way0Dirty_41; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1207 = 7'h2a == reqIndex ? 1'h0 : way0Dirty_42; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1208 = 7'h2b == reqIndex ? 1'h0 : way0Dirty_43; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1209 = 7'h2c == reqIndex ? 1'h0 : way0Dirty_44; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1210 = 7'h2d == reqIndex ? 1'h0 : way0Dirty_45; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1211 = 7'h2e == reqIndex ? 1'h0 : way0Dirty_46; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1212 = 7'h2f == reqIndex ? 1'h0 : way0Dirty_47; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1213 = 7'h30 == reqIndex ? 1'h0 : way0Dirty_48; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1214 = 7'h31 == reqIndex ? 1'h0 : way0Dirty_49; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1215 = 7'h32 == reqIndex ? 1'h0 : way0Dirty_50; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1216 = 7'h33 == reqIndex ? 1'h0 : way0Dirty_51; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1217 = 7'h34 == reqIndex ? 1'h0 : way0Dirty_52; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1218 = 7'h35 == reqIndex ? 1'h0 : way0Dirty_53; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1219 = 7'h36 == reqIndex ? 1'h0 : way0Dirty_54; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1220 = 7'h37 == reqIndex ? 1'h0 : way0Dirty_55; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1221 = 7'h38 == reqIndex ? 1'h0 : way0Dirty_56; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1222 = 7'h39 == reqIndex ? 1'h0 : way0Dirty_57; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1223 = 7'h3a == reqIndex ? 1'h0 : way0Dirty_58; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1224 = 7'h3b == reqIndex ? 1'h0 : way0Dirty_59; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1225 = 7'h3c == reqIndex ? 1'h0 : way0Dirty_60; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1226 = 7'h3d == reqIndex ? 1'h0 : way0Dirty_61; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1227 = 7'h3e == reqIndex ? 1'h0 : way0Dirty_62; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1228 = 7'h3f == reqIndex ? 1'h0 : way0Dirty_63; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1229 = 7'h40 == reqIndex ? 1'h0 : way0Dirty_64; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1230 = 7'h41 == reqIndex ? 1'h0 : way0Dirty_65; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1231 = 7'h42 == reqIndex ? 1'h0 : way0Dirty_66; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1232 = 7'h43 == reqIndex ? 1'h0 : way0Dirty_67; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1233 = 7'h44 == reqIndex ? 1'h0 : way0Dirty_68; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1234 = 7'h45 == reqIndex ? 1'h0 : way0Dirty_69; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1235 = 7'h46 == reqIndex ? 1'h0 : way0Dirty_70; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1236 = 7'h47 == reqIndex ? 1'h0 : way0Dirty_71; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1237 = 7'h48 == reqIndex ? 1'h0 : way0Dirty_72; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1238 = 7'h49 == reqIndex ? 1'h0 : way0Dirty_73; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1239 = 7'h4a == reqIndex ? 1'h0 : way0Dirty_74; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1240 = 7'h4b == reqIndex ? 1'h0 : way0Dirty_75; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1241 = 7'h4c == reqIndex ? 1'h0 : way0Dirty_76; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1242 = 7'h4d == reqIndex ? 1'h0 : way0Dirty_77; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1243 = 7'h4e == reqIndex ? 1'h0 : way0Dirty_78; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1244 = 7'h4f == reqIndex ? 1'h0 : way0Dirty_79; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1245 = 7'h50 == reqIndex ? 1'h0 : way0Dirty_80; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1246 = 7'h51 == reqIndex ? 1'h0 : way0Dirty_81; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1247 = 7'h52 == reqIndex ? 1'h0 : way0Dirty_82; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1248 = 7'h53 == reqIndex ? 1'h0 : way0Dirty_83; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1249 = 7'h54 == reqIndex ? 1'h0 : way0Dirty_84; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1250 = 7'h55 == reqIndex ? 1'h0 : way0Dirty_85; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1251 = 7'h56 == reqIndex ? 1'h0 : way0Dirty_86; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1252 = 7'h57 == reqIndex ? 1'h0 : way0Dirty_87; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1253 = 7'h58 == reqIndex ? 1'h0 : way0Dirty_88; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1254 = 7'h59 == reqIndex ? 1'h0 : way0Dirty_89; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1255 = 7'h5a == reqIndex ? 1'h0 : way0Dirty_90; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1256 = 7'h5b == reqIndex ? 1'h0 : way0Dirty_91; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1257 = 7'h5c == reqIndex ? 1'h0 : way0Dirty_92; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1258 = 7'h5d == reqIndex ? 1'h0 : way0Dirty_93; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1259 = 7'h5e == reqIndex ? 1'h0 : way0Dirty_94; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1260 = 7'h5f == reqIndex ? 1'h0 : way0Dirty_95; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1261 = 7'h60 == reqIndex ? 1'h0 : way0Dirty_96; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1262 = 7'h61 == reqIndex ? 1'h0 : way0Dirty_97; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1263 = 7'h62 == reqIndex ? 1'h0 : way0Dirty_98; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1264 = 7'h63 == reqIndex ? 1'h0 : way0Dirty_99; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1265 = 7'h64 == reqIndex ? 1'h0 : way0Dirty_100; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1266 = 7'h65 == reqIndex ? 1'h0 : way0Dirty_101; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1267 = 7'h66 == reqIndex ? 1'h0 : way0Dirty_102; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1268 = 7'h67 == reqIndex ? 1'h0 : way0Dirty_103; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1269 = 7'h68 == reqIndex ? 1'h0 : way0Dirty_104; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1270 = 7'h69 == reqIndex ? 1'h0 : way0Dirty_105; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1271 = 7'h6a == reqIndex ? 1'h0 : way0Dirty_106; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1272 = 7'h6b == reqIndex ? 1'h0 : way0Dirty_107; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1273 = 7'h6c == reqIndex ? 1'h0 : way0Dirty_108; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1274 = 7'h6d == reqIndex ? 1'h0 : way0Dirty_109; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1275 = 7'h6e == reqIndex ? 1'h0 : way0Dirty_110; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1276 = 7'h6f == reqIndex ? 1'h0 : way0Dirty_111; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1277 = 7'h70 == reqIndex ? 1'h0 : way0Dirty_112; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1278 = 7'h71 == reqIndex ? 1'h0 : way0Dirty_113; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1279 = 7'h72 == reqIndex ? 1'h0 : way0Dirty_114; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1280 = 7'h73 == reqIndex ? 1'h0 : way0Dirty_115; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1281 = 7'h74 == reqIndex ? 1'h0 : way0Dirty_116; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1282 = 7'h75 == reqIndex ? 1'h0 : way0Dirty_117; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1283 = 7'h76 == reqIndex ? 1'h0 : way0Dirty_118; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1284 = 7'h77 == reqIndex ? 1'h0 : way0Dirty_119; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1285 = 7'h78 == reqIndex ? 1'h0 : way0Dirty_120; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1286 = 7'h79 == reqIndex ? 1'h0 : way0Dirty_121; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1287 = 7'h7a == reqIndex ? 1'h0 : way0Dirty_122; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1288 = 7'h7b == reqIndex ? 1'h0 : way0Dirty_123; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1289 = 7'h7c == reqIndex ? 1'h0 : way0Dirty_124; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1290 = 7'h7d == reqIndex ? 1'h0 : way0Dirty_125; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1291 = 7'h7e == reqIndex ? 1'h0 : way0Dirty_126; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1292 = 7'h7f == reqIndex ? 1'h0 : way0Dirty_127; // @[DCache.scala 186:{27,27} 37:26]
  wire  _GEN_1549 = _GEN_4749 | way1Dirty_0; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1550 = _GEN_4750 | way1Dirty_1; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1551 = _GEN_4751 | way1Dirty_2; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1552 = _GEN_4752 | way1Dirty_3; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1553 = _GEN_4753 | way1Dirty_4; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1554 = _GEN_4754 | way1Dirty_5; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1555 = _GEN_4755 | way1Dirty_6; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1556 = _GEN_4756 | way1Dirty_7; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1557 = _GEN_4757 | way1Dirty_8; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1558 = _GEN_4758 | way1Dirty_9; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1559 = _GEN_4759 | way1Dirty_10; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1560 = _GEN_4760 | way1Dirty_11; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1561 = _GEN_4761 | way1Dirty_12; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1562 = _GEN_4762 | way1Dirty_13; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1563 = _GEN_4763 | way1Dirty_14; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1564 = _GEN_4764 | way1Dirty_15; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1565 = _GEN_4765 | way1Dirty_16; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1566 = _GEN_4766 | way1Dirty_17; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1567 = _GEN_4767 | way1Dirty_18; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1568 = _GEN_4768 | way1Dirty_19; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1569 = _GEN_4769 | way1Dirty_20; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1570 = _GEN_4770 | way1Dirty_21; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1571 = _GEN_4771 | way1Dirty_22; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1572 = _GEN_4772 | way1Dirty_23; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1573 = _GEN_4773 | way1Dirty_24; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1574 = _GEN_4774 | way1Dirty_25; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1575 = _GEN_4775 | way1Dirty_26; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1576 = _GEN_4776 | way1Dirty_27; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1577 = _GEN_4777 | way1Dirty_28; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1578 = _GEN_4778 | way1Dirty_29; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1579 = _GEN_4779 | way1Dirty_30; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1580 = _GEN_4780 | way1Dirty_31; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1581 = _GEN_4781 | way1Dirty_32; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1582 = _GEN_4782 | way1Dirty_33; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1583 = _GEN_4783 | way1Dirty_34; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1584 = _GEN_4784 | way1Dirty_35; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1585 = _GEN_4785 | way1Dirty_36; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1586 = _GEN_4786 | way1Dirty_37; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1587 = _GEN_4787 | way1Dirty_38; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1588 = _GEN_4788 | way1Dirty_39; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1589 = _GEN_4789 | way1Dirty_40; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1590 = _GEN_4790 | way1Dirty_41; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1591 = _GEN_4791 | way1Dirty_42; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1592 = _GEN_4792 | way1Dirty_43; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1593 = _GEN_4793 | way1Dirty_44; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1594 = _GEN_4794 | way1Dirty_45; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1595 = _GEN_4795 | way1Dirty_46; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1596 = _GEN_4796 | way1Dirty_47; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1597 = _GEN_4797 | way1Dirty_48; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1598 = _GEN_4798 | way1Dirty_49; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1599 = _GEN_4799 | way1Dirty_50; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1600 = _GEN_4800 | way1Dirty_51; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1601 = _GEN_4801 | way1Dirty_52; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1602 = _GEN_4802 | way1Dirty_53; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1603 = _GEN_4803 | way1Dirty_54; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1604 = _GEN_4804 | way1Dirty_55; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1605 = _GEN_4805 | way1Dirty_56; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1606 = _GEN_4806 | way1Dirty_57; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1607 = _GEN_4807 | way1Dirty_58; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1608 = _GEN_4808 | way1Dirty_59; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1609 = _GEN_4809 | way1Dirty_60; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1610 = _GEN_4810 | way1Dirty_61; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1611 = _GEN_4811 | way1Dirty_62; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1612 = _GEN_4812 | way1Dirty_63; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1613 = _GEN_4813 | way1Dirty_64; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1614 = _GEN_4814 | way1Dirty_65; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1615 = _GEN_4815 | way1Dirty_66; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1616 = _GEN_4816 | way1Dirty_67; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1617 = _GEN_4817 | way1Dirty_68; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1618 = _GEN_4818 | way1Dirty_69; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1619 = _GEN_4819 | way1Dirty_70; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1620 = _GEN_4820 | way1Dirty_71; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1621 = _GEN_4821 | way1Dirty_72; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1622 = _GEN_4822 | way1Dirty_73; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1623 = _GEN_4823 | way1Dirty_74; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1624 = _GEN_4824 | way1Dirty_75; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1625 = _GEN_4825 | way1Dirty_76; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1626 = _GEN_4826 | way1Dirty_77; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1627 = _GEN_4827 | way1Dirty_78; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1628 = _GEN_4828 | way1Dirty_79; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1629 = _GEN_4829 | way1Dirty_80; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1630 = _GEN_4830 | way1Dirty_81; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1631 = _GEN_4831 | way1Dirty_82; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1632 = _GEN_4832 | way1Dirty_83; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1633 = _GEN_4833 | way1Dirty_84; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1634 = _GEN_4834 | way1Dirty_85; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1635 = _GEN_4835 | way1Dirty_86; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1636 = _GEN_4836 | way1Dirty_87; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1637 = _GEN_4837 | way1Dirty_88; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1638 = _GEN_4838 | way1Dirty_89; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1639 = _GEN_4839 | way1Dirty_90; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1640 = _GEN_4840 | way1Dirty_91; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1641 = _GEN_4841 | way1Dirty_92; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1642 = _GEN_4842 | way1Dirty_93; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1643 = _GEN_4843 | way1Dirty_94; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1644 = _GEN_4844 | way1Dirty_95; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1645 = _GEN_4845 | way1Dirty_96; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1646 = _GEN_4846 | way1Dirty_97; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1647 = _GEN_4847 | way1Dirty_98; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1648 = _GEN_4848 | way1Dirty_99; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1649 = _GEN_4849 | way1Dirty_100; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1650 = _GEN_4850 | way1Dirty_101; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1651 = _GEN_4851 | way1Dirty_102; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1652 = _GEN_4852 | way1Dirty_103; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1653 = _GEN_4853 | way1Dirty_104; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1654 = _GEN_4854 | way1Dirty_105; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1655 = _GEN_4855 | way1Dirty_106; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1656 = _GEN_4856 | way1Dirty_107; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1657 = _GEN_4857 | way1Dirty_108; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1658 = _GEN_4858 | way1Dirty_109; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1659 = _GEN_4859 | way1Dirty_110; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1660 = _GEN_4860 | way1Dirty_111; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1661 = _GEN_4861 | way1Dirty_112; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1662 = _GEN_4862 | way1Dirty_113; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1663 = _GEN_4863 | way1Dirty_114; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1664 = _GEN_4864 | way1Dirty_115; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1665 = _GEN_4865 | way1Dirty_116; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1666 = _GEN_4866 | way1Dirty_117; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1667 = _GEN_4867 | way1Dirty_118; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1668 = _GEN_4868 | way1Dirty_119; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1669 = _GEN_4869 | way1Dirty_120; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1670 = _GEN_4870 | way1Dirty_121; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1671 = _GEN_4871 | way1Dirty_122; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1672 = _GEN_4872 | way1Dirty_123; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1673 = _GEN_4873 | way1Dirty_124; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1674 = _GEN_4874 | way1Dirty_125; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1675 = _GEN_4875 | way1Dirty_126; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1676 = _GEN_4876 | way1Dirty_127; // @[DCache.scala 190:{27,27} 43:26]
  wire  _GEN_1677 = 7'h0 == reqIndex ? 1'h0 : way1Dirty_0; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1678 = 7'h1 == reqIndex ? 1'h0 : way1Dirty_1; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1679 = 7'h2 == reqIndex ? 1'h0 : way1Dirty_2; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1680 = 7'h3 == reqIndex ? 1'h0 : way1Dirty_3; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1681 = 7'h4 == reqIndex ? 1'h0 : way1Dirty_4; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1682 = 7'h5 == reqIndex ? 1'h0 : way1Dirty_5; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1683 = 7'h6 == reqIndex ? 1'h0 : way1Dirty_6; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1684 = 7'h7 == reqIndex ? 1'h0 : way1Dirty_7; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1685 = 7'h8 == reqIndex ? 1'h0 : way1Dirty_8; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1686 = 7'h9 == reqIndex ? 1'h0 : way1Dirty_9; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1687 = 7'ha == reqIndex ? 1'h0 : way1Dirty_10; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1688 = 7'hb == reqIndex ? 1'h0 : way1Dirty_11; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1689 = 7'hc == reqIndex ? 1'h0 : way1Dirty_12; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1690 = 7'hd == reqIndex ? 1'h0 : way1Dirty_13; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1691 = 7'he == reqIndex ? 1'h0 : way1Dirty_14; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1692 = 7'hf == reqIndex ? 1'h0 : way1Dirty_15; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1693 = 7'h10 == reqIndex ? 1'h0 : way1Dirty_16; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1694 = 7'h11 == reqIndex ? 1'h0 : way1Dirty_17; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1695 = 7'h12 == reqIndex ? 1'h0 : way1Dirty_18; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1696 = 7'h13 == reqIndex ? 1'h0 : way1Dirty_19; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1697 = 7'h14 == reqIndex ? 1'h0 : way1Dirty_20; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1698 = 7'h15 == reqIndex ? 1'h0 : way1Dirty_21; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1699 = 7'h16 == reqIndex ? 1'h0 : way1Dirty_22; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1700 = 7'h17 == reqIndex ? 1'h0 : way1Dirty_23; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1701 = 7'h18 == reqIndex ? 1'h0 : way1Dirty_24; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1702 = 7'h19 == reqIndex ? 1'h0 : way1Dirty_25; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1703 = 7'h1a == reqIndex ? 1'h0 : way1Dirty_26; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1704 = 7'h1b == reqIndex ? 1'h0 : way1Dirty_27; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1705 = 7'h1c == reqIndex ? 1'h0 : way1Dirty_28; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1706 = 7'h1d == reqIndex ? 1'h0 : way1Dirty_29; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1707 = 7'h1e == reqIndex ? 1'h0 : way1Dirty_30; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1708 = 7'h1f == reqIndex ? 1'h0 : way1Dirty_31; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1709 = 7'h20 == reqIndex ? 1'h0 : way1Dirty_32; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1710 = 7'h21 == reqIndex ? 1'h0 : way1Dirty_33; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1711 = 7'h22 == reqIndex ? 1'h0 : way1Dirty_34; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1712 = 7'h23 == reqIndex ? 1'h0 : way1Dirty_35; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1713 = 7'h24 == reqIndex ? 1'h0 : way1Dirty_36; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1714 = 7'h25 == reqIndex ? 1'h0 : way1Dirty_37; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1715 = 7'h26 == reqIndex ? 1'h0 : way1Dirty_38; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1716 = 7'h27 == reqIndex ? 1'h0 : way1Dirty_39; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1717 = 7'h28 == reqIndex ? 1'h0 : way1Dirty_40; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1718 = 7'h29 == reqIndex ? 1'h0 : way1Dirty_41; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1719 = 7'h2a == reqIndex ? 1'h0 : way1Dirty_42; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1720 = 7'h2b == reqIndex ? 1'h0 : way1Dirty_43; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1721 = 7'h2c == reqIndex ? 1'h0 : way1Dirty_44; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1722 = 7'h2d == reqIndex ? 1'h0 : way1Dirty_45; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1723 = 7'h2e == reqIndex ? 1'h0 : way1Dirty_46; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1724 = 7'h2f == reqIndex ? 1'h0 : way1Dirty_47; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1725 = 7'h30 == reqIndex ? 1'h0 : way1Dirty_48; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1726 = 7'h31 == reqIndex ? 1'h0 : way1Dirty_49; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1727 = 7'h32 == reqIndex ? 1'h0 : way1Dirty_50; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1728 = 7'h33 == reqIndex ? 1'h0 : way1Dirty_51; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1729 = 7'h34 == reqIndex ? 1'h0 : way1Dirty_52; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1730 = 7'h35 == reqIndex ? 1'h0 : way1Dirty_53; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1731 = 7'h36 == reqIndex ? 1'h0 : way1Dirty_54; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1732 = 7'h37 == reqIndex ? 1'h0 : way1Dirty_55; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1733 = 7'h38 == reqIndex ? 1'h0 : way1Dirty_56; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1734 = 7'h39 == reqIndex ? 1'h0 : way1Dirty_57; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1735 = 7'h3a == reqIndex ? 1'h0 : way1Dirty_58; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1736 = 7'h3b == reqIndex ? 1'h0 : way1Dirty_59; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1737 = 7'h3c == reqIndex ? 1'h0 : way1Dirty_60; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1738 = 7'h3d == reqIndex ? 1'h0 : way1Dirty_61; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1739 = 7'h3e == reqIndex ? 1'h0 : way1Dirty_62; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1740 = 7'h3f == reqIndex ? 1'h0 : way1Dirty_63; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1741 = 7'h40 == reqIndex ? 1'h0 : way1Dirty_64; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1742 = 7'h41 == reqIndex ? 1'h0 : way1Dirty_65; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1743 = 7'h42 == reqIndex ? 1'h0 : way1Dirty_66; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1744 = 7'h43 == reqIndex ? 1'h0 : way1Dirty_67; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1745 = 7'h44 == reqIndex ? 1'h0 : way1Dirty_68; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1746 = 7'h45 == reqIndex ? 1'h0 : way1Dirty_69; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1747 = 7'h46 == reqIndex ? 1'h0 : way1Dirty_70; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1748 = 7'h47 == reqIndex ? 1'h0 : way1Dirty_71; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1749 = 7'h48 == reqIndex ? 1'h0 : way1Dirty_72; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1750 = 7'h49 == reqIndex ? 1'h0 : way1Dirty_73; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1751 = 7'h4a == reqIndex ? 1'h0 : way1Dirty_74; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1752 = 7'h4b == reqIndex ? 1'h0 : way1Dirty_75; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1753 = 7'h4c == reqIndex ? 1'h0 : way1Dirty_76; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1754 = 7'h4d == reqIndex ? 1'h0 : way1Dirty_77; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1755 = 7'h4e == reqIndex ? 1'h0 : way1Dirty_78; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1756 = 7'h4f == reqIndex ? 1'h0 : way1Dirty_79; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1757 = 7'h50 == reqIndex ? 1'h0 : way1Dirty_80; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1758 = 7'h51 == reqIndex ? 1'h0 : way1Dirty_81; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1759 = 7'h52 == reqIndex ? 1'h0 : way1Dirty_82; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1760 = 7'h53 == reqIndex ? 1'h0 : way1Dirty_83; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1761 = 7'h54 == reqIndex ? 1'h0 : way1Dirty_84; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1762 = 7'h55 == reqIndex ? 1'h0 : way1Dirty_85; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1763 = 7'h56 == reqIndex ? 1'h0 : way1Dirty_86; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1764 = 7'h57 == reqIndex ? 1'h0 : way1Dirty_87; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1765 = 7'h58 == reqIndex ? 1'h0 : way1Dirty_88; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1766 = 7'h59 == reqIndex ? 1'h0 : way1Dirty_89; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1767 = 7'h5a == reqIndex ? 1'h0 : way1Dirty_90; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1768 = 7'h5b == reqIndex ? 1'h0 : way1Dirty_91; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1769 = 7'h5c == reqIndex ? 1'h0 : way1Dirty_92; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1770 = 7'h5d == reqIndex ? 1'h0 : way1Dirty_93; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1771 = 7'h5e == reqIndex ? 1'h0 : way1Dirty_94; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1772 = 7'h5f == reqIndex ? 1'h0 : way1Dirty_95; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1773 = 7'h60 == reqIndex ? 1'h0 : way1Dirty_96; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1774 = 7'h61 == reqIndex ? 1'h0 : way1Dirty_97; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1775 = 7'h62 == reqIndex ? 1'h0 : way1Dirty_98; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1776 = 7'h63 == reqIndex ? 1'h0 : way1Dirty_99; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1777 = 7'h64 == reqIndex ? 1'h0 : way1Dirty_100; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1778 = 7'h65 == reqIndex ? 1'h0 : way1Dirty_101; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1779 = 7'h66 == reqIndex ? 1'h0 : way1Dirty_102; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1780 = 7'h67 == reqIndex ? 1'h0 : way1Dirty_103; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1781 = 7'h68 == reqIndex ? 1'h0 : way1Dirty_104; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1782 = 7'h69 == reqIndex ? 1'h0 : way1Dirty_105; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1783 = 7'h6a == reqIndex ? 1'h0 : way1Dirty_106; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1784 = 7'h6b == reqIndex ? 1'h0 : way1Dirty_107; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1785 = 7'h6c == reqIndex ? 1'h0 : way1Dirty_108; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1786 = 7'h6d == reqIndex ? 1'h0 : way1Dirty_109; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1787 = 7'h6e == reqIndex ? 1'h0 : way1Dirty_110; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1788 = 7'h6f == reqIndex ? 1'h0 : way1Dirty_111; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1789 = 7'h70 == reqIndex ? 1'h0 : way1Dirty_112; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1790 = 7'h71 == reqIndex ? 1'h0 : way1Dirty_113; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1791 = 7'h72 == reqIndex ? 1'h0 : way1Dirty_114; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1792 = 7'h73 == reqIndex ? 1'h0 : way1Dirty_115; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1793 = 7'h74 == reqIndex ? 1'h0 : way1Dirty_116; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1794 = 7'h75 == reqIndex ? 1'h0 : way1Dirty_117; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1795 = 7'h76 == reqIndex ? 1'h0 : way1Dirty_118; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1796 = 7'h77 == reqIndex ? 1'h0 : way1Dirty_119; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1797 = 7'h78 == reqIndex ? 1'h0 : way1Dirty_120; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1798 = 7'h79 == reqIndex ? 1'h0 : way1Dirty_121; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1799 = 7'h7a == reqIndex ? 1'h0 : way1Dirty_122; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1800 = 7'h7b == reqIndex ? 1'h0 : way1Dirty_123; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1801 = 7'h7c == reqIndex ? 1'h0 : way1Dirty_124; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1802 = 7'h7d == reqIndex ? 1'h0 : way1Dirty_125; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1803 = 7'h7e == reqIndex ? 1'h0 : way1Dirty_126; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1804 = 7'h7f == reqIndex ? 1'h0 : way1Dirty_127; // @[DCache.scala 192:{27,27} 43:26]
  wire  _GEN_1805 = _T_10 ? _GEN_1677 : way1Dirty_0; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1806 = _T_10 ? _GEN_1678 : way1Dirty_1; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1807 = _T_10 ? _GEN_1679 : way1Dirty_2; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1808 = _T_10 ? _GEN_1680 : way1Dirty_3; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1809 = _T_10 ? _GEN_1681 : way1Dirty_4; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1810 = _T_10 ? _GEN_1682 : way1Dirty_5; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1811 = _T_10 ? _GEN_1683 : way1Dirty_6; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1812 = _T_10 ? _GEN_1684 : way1Dirty_7; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1813 = _T_10 ? _GEN_1685 : way1Dirty_8; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1814 = _T_10 ? _GEN_1686 : way1Dirty_9; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1815 = _T_10 ? _GEN_1687 : way1Dirty_10; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1816 = _T_10 ? _GEN_1688 : way1Dirty_11; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1817 = _T_10 ? _GEN_1689 : way1Dirty_12; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1818 = _T_10 ? _GEN_1690 : way1Dirty_13; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1819 = _T_10 ? _GEN_1691 : way1Dirty_14; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1820 = _T_10 ? _GEN_1692 : way1Dirty_15; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1821 = _T_10 ? _GEN_1693 : way1Dirty_16; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1822 = _T_10 ? _GEN_1694 : way1Dirty_17; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1823 = _T_10 ? _GEN_1695 : way1Dirty_18; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1824 = _T_10 ? _GEN_1696 : way1Dirty_19; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1825 = _T_10 ? _GEN_1697 : way1Dirty_20; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1826 = _T_10 ? _GEN_1698 : way1Dirty_21; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1827 = _T_10 ? _GEN_1699 : way1Dirty_22; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1828 = _T_10 ? _GEN_1700 : way1Dirty_23; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1829 = _T_10 ? _GEN_1701 : way1Dirty_24; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1830 = _T_10 ? _GEN_1702 : way1Dirty_25; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1831 = _T_10 ? _GEN_1703 : way1Dirty_26; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1832 = _T_10 ? _GEN_1704 : way1Dirty_27; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1833 = _T_10 ? _GEN_1705 : way1Dirty_28; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1834 = _T_10 ? _GEN_1706 : way1Dirty_29; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1835 = _T_10 ? _GEN_1707 : way1Dirty_30; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1836 = _T_10 ? _GEN_1708 : way1Dirty_31; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1837 = _T_10 ? _GEN_1709 : way1Dirty_32; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1838 = _T_10 ? _GEN_1710 : way1Dirty_33; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1839 = _T_10 ? _GEN_1711 : way1Dirty_34; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1840 = _T_10 ? _GEN_1712 : way1Dirty_35; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1841 = _T_10 ? _GEN_1713 : way1Dirty_36; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1842 = _T_10 ? _GEN_1714 : way1Dirty_37; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1843 = _T_10 ? _GEN_1715 : way1Dirty_38; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1844 = _T_10 ? _GEN_1716 : way1Dirty_39; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1845 = _T_10 ? _GEN_1717 : way1Dirty_40; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1846 = _T_10 ? _GEN_1718 : way1Dirty_41; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1847 = _T_10 ? _GEN_1719 : way1Dirty_42; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1848 = _T_10 ? _GEN_1720 : way1Dirty_43; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1849 = _T_10 ? _GEN_1721 : way1Dirty_44; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1850 = _T_10 ? _GEN_1722 : way1Dirty_45; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1851 = _T_10 ? _GEN_1723 : way1Dirty_46; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1852 = _T_10 ? _GEN_1724 : way1Dirty_47; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1853 = _T_10 ? _GEN_1725 : way1Dirty_48; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1854 = _T_10 ? _GEN_1726 : way1Dirty_49; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1855 = _T_10 ? _GEN_1727 : way1Dirty_50; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1856 = _T_10 ? _GEN_1728 : way1Dirty_51; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1857 = _T_10 ? _GEN_1729 : way1Dirty_52; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1858 = _T_10 ? _GEN_1730 : way1Dirty_53; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1859 = _T_10 ? _GEN_1731 : way1Dirty_54; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1860 = _T_10 ? _GEN_1732 : way1Dirty_55; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1861 = _T_10 ? _GEN_1733 : way1Dirty_56; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1862 = _T_10 ? _GEN_1734 : way1Dirty_57; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1863 = _T_10 ? _GEN_1735 : way1Dirty_58; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1864 = _T_10 ? _GEN_1736 : way1Dirty_59; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1865 = _T_10 ? _GEN_1737 : way1Dirty_60; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1866 = _T_10 ? _GEN_1738 : way1Dirty_61; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1867 = _T_10 ? _GEN_1739 : way1Dirty_62; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1868 = _T_10 ? _GEN_1740 : way1Dirty_63; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1869 = _T_10 ? _GEN_1741 : way1Dirty_64; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1870 = _T_10 ? _GEN_1742 : way1Dirty_65; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1871 = _T_10 ? _GEN_1743 : way1Dirty_66; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1872 = _T_10 ? _GEN_1744 : way1Dirty_67; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1873 = _T_10 ? _GEN_1745 : way1Dirty_68; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1874 = _T_10 ? _GEN_1746 : way1Dirty_69; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1875 = _T_10 ? _GEN_1747 : way1Dirty_70; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1876 = _T_10 ? _GEN_1748 : way1Dirty_71; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1877 = _T_10 ? _GEN_1749 : way1Dirty_72; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1878 = _T_10 ? _GEN_1750 : way1Dirty_73; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1879 = _T_10 ? _GEN_1751 : way1Dirty_74; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1880 = _T_10 ? _GEN_1752 : way1Dirty_75; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1881 = _T_10 ? _GEN_1753 : way1Dirty_76; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1882 = _T_10 ? _GEN_1754 : way1Dirty_77; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1883 = _T_10 ? _GEN_1755 : way1Dirty_78; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1884 = _T_10 ? _GEN_1756 : way1Dirty_79; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1885 = _T_10 ? _GEN_1757 : way1Dirty_80; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1886 = _T_10 ? _GEN_1758 : way1Dirty_81; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1887 = _T_10 ? _GEN_1759 : way1Dirty_82; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1888 = _T_10 ? _GEN_1760 : way1Dirty_83; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1889 = _T_10 ? _GEN_1761 : way1Dirty_84; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1890 = _T_10 ? _GEN_1762 : way1Dirty_85; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1891 = _T_10 ? _GEN_1763 : way1Dirty_86; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1892 = _T_10 ? _GEN_1764 : way1Dirty_87; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1893 = _T_10 ? _GEN_1765 : way1Dirty_88; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1894 = _T_10 ? _GEN_1766 : way1Dirty_89; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1895 = _T_10 ? _GEN_1767 : way1Dirty_90; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1896 = _T_10 ? _GEN_1768 : way1Dirty_91; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1897 = _T_10 ? _GEN_1769 : way1Dirty_92; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1898 = _T_10 ? _GEN_1770 : way1Dirty_93; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1899 = _T_10 ? _GEN_1771 : way1Dirty_94; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1900 = _T_10 ? _GEN_1772 : way1Dirty_95; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1901 = _T_10 ? _GEN_1773 : way1Dirty_96; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1902 = _T_10 ? _GEN_1774 : way1Dirty_97; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1903 = _T_10 ? _GEN_1775 : way1Dirty_98; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1904 = _T_10 ? _GEN_1776 : way1Dirty_99; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1905 = _T_10 ? _GEN_1777 : way1Dirty_100; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1906 = _T_10 ? _GEN_1778 : way1Dirty_101; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1907 = _T_10 ? _GEN_1779 : way1Dirty_102; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1908 = _T_10 ? _GEN_1780 : way1Dirty_103; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1909 = _T_10 ? _GEN_1781 : way1Dirty_104; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1910 = _T_10 ? _GEN_1782 : way1Dirty_105; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1911 = _T_10 ? _GEN_1783 : way1Dirty_106; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1912 = _T_10 ? _GEN_1784 : way1Dirty_107; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1913 = _T_10 ? _GEN_1785 : way1Dirty_108; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1914 = _T_10 ? _GEN_1786 : way1Dirty_109; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1915 = _T_10 ? _GEN_1787 : way1Dirty_110; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1916 = _T_10 ? _GEN_1788 : way1Dirty_111; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1917 = _T_10 ? _GEN_1789 : way1Dirty_112; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1918 = _T_10 ? _GEN_1790 : way1Dirty_113; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1919 = _T_10 ? _GEN_1791 : way1Dirty_114; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1920 = _T_10 ? _GEN_1792 : way1Dirty_115; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1921 = _T_10 ? _GEN_1793 : way1Dirty_116; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1922 = _T_10 ? _GEN_1794 : way1Dirty_117; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1923 = _T_10 ? _GEN_1795 : way1Dirty_118; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1924 = _T_10 ? _GEN_1796 : way1Dirty_119; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1925 = _T_10 ? _GEN_1797 : way1Dirty_120; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1926 = _T_10 ? _GEN_1798 : way1Dirty_121; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1927 = _T_10 ? _GEN_1799 : way1Dirty_122; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1928 = _T_10 ? _GEN_1800 : way1Dirty_123; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1929 = _T_10 ? _GEN_1801 : way1Dirty_124; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1930 = _T_10 ? _GEN_1802 : way1Dirty_125; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1931 = _T_10 ? _GEN_1803 : way1Dirty_126; // @[DCache.scala 191:45 43:26]
  wire  _GEN_1932 = _T_10 ? _GEN_1804 : way1Dirty_127; // @[DCache.scala 191:45 43:26]
  wire  sDoneEn = state == 3'h6; // @[DCache.scala 196:23]
  wire  _GEN_2445 = _GEN_4749 | way0V_0; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2446 = _GEN_4750 | way0V_1; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2447 = _GEN_4751 | way0V_2; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2448 = _GEN_4752 | way0V_3; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2449 = _GEN_4753 | way0V_4; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2450 = _GEN_4754 | way0V_5; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2451 = _GEN_4755 | way0V_6; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2452 = _GEN_4756 | way0V_7; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2453 = _GEN_4757 | way0V_8; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2454 = _GEN_4758 | way0V_9; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2455 = _GEN_4759 | way0V_10; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2456 = _GEN_4760 | way0V_11; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2457 = _GEN_4761 | way0V_12; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2458 = _GEN_4762 | way0V_13; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2459 = _GEN_4763 | way0V_14; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2460 = _GEN_4764 | way0V_15; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2461 = _GEN_4765 | way0V_16; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2462 = _GEN_4766 | way0V_17; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2463 = _GEN_4767 | way0V_18; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2464 = _GEN_4768 | way0V_19; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2465 = _GEN_4769 | way0V_20; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2466 = _GEN_4770 | way0V_21; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2467 = _GEN_4771 | way0V_22; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2468 = _GEN_4772 | way0V_23; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2469 = _GEN_4773 | way0V_24; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2470 = _GEN_4774 | way0V_25; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2471 = _GEN_4775 | way0V_26; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2472 = _GEN_4776 | way0V_27; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2473 = _GEN_4777 | way0V_28; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2474 = _GEN_4778 | way0V_29; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2475 = _GEN_4779 | way0V_30; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2476 = _GEN_4780 | way0V_31; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2477 = _GEN_4781 | way0V_32; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2478 = _GEN_4782 | way0V_33; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2479 = _GEN_4783 | way0V_34; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2480 = _GEN_4784 | way0V_35; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2481 = _GEN_4785 | way0V_36; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2482 = _GEN_4786 | way0V_37; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2483 = _GEN_4787 | way0V_38; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2484 = _GEN_4788 | way0V_39; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2485 = _GEN_4789 | way0V_40; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2486 = _GEN_4790 | way0V_41; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2487 = _GEN_4791 | way0V_42; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2488 = _GEN_4792 | way0V_43; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2489 = _GEN_4793 | way0V_44; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2490 = _GEN_4794 | way0V_45; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2491 = _GEN_4795 | way0V_46; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2492 = _GEN_4796 | way0V_47; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2493 = _GEN_4797 | way0V_48; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2494 = _GEN_4798 | way0V_49; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2495 = _GEN_4799 | way0V_50; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2496 = _GEN_4800 | way0V_51; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2497 = _GEN_4801 | way0V_52; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2498 = _GEN_4802 | way0V_53; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2499 = _GEN_4803 | way0V_54; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2500 = _GEN_4804 | way0V_55; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2501 = _GEN_4805 | way0V_56; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2502 = _GEN_4806 | way0V_57; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2503 = _GEN_4807 | way0V_58; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2504 = _GEN_4808 | way0V_59; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2505 = _GEN_4809 | way0V_60; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2506 = _GEN_4810 | way0V_61; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2507 = _GEN_4811 | way0V_62; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2508 = _GEN_4812 | way0V_63; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2509 = _GEN_4813 | way0V_64; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2510 = _GEN_4814 | way0V_65; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2511 = _GEN_4815 | way0V_66; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2512 = _GEN_4816 | way0V_67; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2513 = _GEN_4817 | way0V_68; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2514 = _GEN_4818 | way0V_69; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2515 = _GEN_4819 | way0V_70; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2516 = _GEN_4820 | way0V_71; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2517 = _GEN_4821 | way0V_72; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2518 = _GEN_4822 | way0V_73; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2519 = _GEN_4823 | way0V_74; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2520 = _GEN_4824 | way0V_75; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2521 = _GEN_4825 | way0V_76; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2522 = _GEN_4826 | way0V_77; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2523 = _GEN_4827 | way0V_78; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2524 = _GEN_4828 | way0V_79; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2525 = _GEN_4829 | way0V_80; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2526 = _GEN_4830 | way0V_81; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2527 = _GEN_4831 | way0V_82; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2528 = _GEN_4832 | way0V_83; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2529 = _GEN_4833 | way0V_84; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2530 = _GEN_4834 | way0V_85; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2531 = _GEN_4835 | way0V_86; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2532 = _GEN_4836 | way0V_87; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2533 = _GEN_4837 | way0V_88; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2534 = _GEN_4838 | way0V_89; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2535 = _GEN_4839 | way0V_90; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2536 = _GEN_4840 | way0V_91; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2537 = _GEN_4841 | way0V_92; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2538 = _GEN_4842 | way0V_93; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2539 = _GEN_4843 | way0V_94; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2540 = _GEN_4844 | way0V_95; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2541 = _GEN_4845 | way0V_96; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2542 = _GEN_4846 | way0V_97; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2543 = _GEN_4847 | way0V_98; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2544 = _GEN_4848 | way0V_99; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2545 = _GEN_4849 | way0V_100; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2546 = _GEN_4850 | way0V_101; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2547 = _GEN_4851 | way0V_102; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2548 = _GEN_4852 | way0V_103; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2549 = _GEN_4853 | way0V_104; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2550 = _GEN_4854 | way0V_105; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2551 = _GEN_4855 | way0V_106; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2552 = _GEN_4856 | way0V_107; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2553 = _GEN_4857 | way0V_108; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2554 = _GEN_4858 | way0V_109; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2555 = _GEN_4859 | way0V_110; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2556 = _GEN_4860 | way0V_111; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2557 = _GEN_4861 | way0V_112; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2558 = _GEN_4862 | way0V_113; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2559 = _GEN_4863 | way0V_114; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2560 = _GEN_4864 | way0V_115; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2561 = _GEN_4865 | way0V_116; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2562 = _GEN_4866 | way0V_117; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2563 = _GEN_4867 | way0V_118; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2564 = _GEN_4868 | way0V_119; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2565 = _GEN_4869 | way0V_120; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2566 = _GEN_4870 | way0V_121; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2567 = _GEN_4871 | way0V_122; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2568 = _GEN_4872 | way0V_123; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2569 = _GEN_4873 | way0V_124; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2570 = _GEN_4874 | way0V_125; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2571 = _GEN_4875 | way0V_126; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2572 = _GEN_4876 | way0V_127; // @[DCache.scala 199:{21,21} 33:26]
  wire  _GEN_2701 = _GEN_4749 | way0Age_0; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2702 = _GEN_4750 | way0Age_1; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2703 = _GEN_4751 | way0Age_2; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2704 = _GEN_4752 | way0Age_3; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2705 = _GEN_4753 | way0Age_4; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2706 = _GEN_4754 | way0Age_5; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2707 = _GEN_4755 | way0Age_6; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2708 = _GEN_4756 | way0Age_7; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2709 = _GEN_4757 | way0Age_8; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2710 = _GEN_4758 | way0Age_9; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2711 = _GEN_4759 | way0Age_10; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2712 = _GEN_4760 | way0Age_11; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2713 = _GEN_4761 | way0Age_12; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2714 = _GEN_4762 | way0Age_13; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2715 = _GEN_4763 | way0Age_14; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2716 = _GEN_4764 | way0Age_15; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2717 = _GEN_4765 | way0Age_16; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2718 = _GEN_4766 | way0Age_17; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2719 = _GEN_4767 | way0Age_18; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2720 = _GEN_4768 | way0Age_19; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2721 = _GEN_4769 | way0Age_20; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2722 = _GEN_4770 | way0Age_21; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2723 = _GEN_4771 | way0Age_22; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2724 = _GEN_4772 | way0Age_23; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2725 = _GEN_4773 | way0Age_24; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2726 = _GEN_4774 | way0Age_25; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2727 = _GEN_4775 | way0Age_26; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2728 = _GEN_4776 | way0Age_27; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2729 = _GEN_4777 | way0Age_28; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2730 = _GEN_4778 | way0Age_29; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2731 = _GEN_4779 | way0Age_30; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2732 = _GEN_4780 | way0Age_31; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2733 = _GEN_4781 | way0Age_32; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2734 = _GEN_4782 | way0Age_33; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2735 = _GEN_4783 | way0Age_34; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2736 = _GEN_4784 | way0Age_35; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2737 = _GEN_4785 | way0Age_36; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2738 = _GEN_4786 | way0Age_37; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2739 = _GEN_4787 | way0Age_38; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2740 = _GEN_4788 | way0Age_39; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2741 = _GEN_4789 | way0Age_40; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2742 = _GEN_4790 | way0Age_41; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2743 = _GEN_4791 | way0Age_42; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2744 = _GEN_4792 | way0Age_43; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2745 = _GEN_4793 | way0Age_44; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2746 = _GEN_4794 | way0Age_45; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2747 = _GEN_4795 | way0Age_46; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2748 = _GEN_4796 | way0Age_47; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2749 = _GEN_4797 | way0Age_48; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2750 = _GEN_4798 | way0Age_49; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2751 = _GEN_4799 | way0Age_50; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2752 = _GEN_4800 | way0Age_51; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2753 = _GEN_4801 | way0Age_52; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2754 = _GEN_4802 | way0Age_53; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2755 = _GEN_4803 | way0Age_54; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2756 = _GEN_4804 | way0Age_55; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2757 = _GEN_4805 | way0Age_56; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2758 = _GEN_4806 | way0Age_57; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2759 = _GEN_4807 | way0Age_58; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2760 = _GEN_4808 | way0Age_59; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2761 = _GEN_4809 | way0Age_60; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2762 = _GEN_4810 | way0Age_61; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2763 = _GEN_4811 | way0Age_62; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2764 = _GEN_4812 | way0Age_63; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2765 = _GEN_4813 | way0Age_64; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2766 = _GEN_4814 | way0Age_65; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2767 = _GEN_4815 | way0Age_66; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2768 = _GEN_4816 | way0Age_67; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2769 = _GEN_4817 | way0Age_68; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2770 = _GEN_4818 | way0Age_69; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2771 = _GEN_4819 | way0Age_70; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2772 = _GEN_4820 | way0Age_71; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2773 = _GEN_4821 | way0Age_72; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2774 = _GEN_4822 | way0Age_73; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2775 = _GEN_4823 | way0Age_74; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2776 = _GEN_4824 | way0Age_75; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2777 = _GEN_4825 | way0Age_76; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2778 = _GEN_4826 | way0Age_77; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2779 = _GEN_4827 | way0Age_78; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2780 = _GEN_4828 | way0Age_79; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2781 = _GEN_4829 | way0Age_80; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2782 = _GEN_4830 | way0Age_81; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2783 = _GEN_4831 | way0Age_82; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2784 = _GEN_4832 | way0Age_83; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2785 = _GEN_4833 | way0Age_84; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2786 = _GEN_4834 | way0Age_85; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2787 = _GEN_4835 | way0Age_86; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2788 = _GEN_4836 | way0Age_87; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2789 = _GEN_4837 | way0Age_88; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2790 = _GEN_4838 | way0Age_89; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2791 = _GEN_4839 | way0Age_90; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2792 = _GEN_4840 | way0Age_91; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2793 = _GEN_4841 | way0Age_92; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2794 = _GEN_4842 | way0Age_93; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2795 = _GEN_4843 | way0Age_94; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2796 = _GEN_4844 | way0Age_95; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2797 = _GEN_4845 | way0Age_96; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2798 = _GEN_4846 | way0Age_97; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2799 = _GEN_4847 | way0Age_98; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2800 = _GEN_4848 | way0Age_99; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2801 = _GEN_4849 | way0Age_100; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2802 = _GEN_4850 | way0Age_101; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2803 = _GEN_4851 | way0Age_102; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2804 = _GEN_4852 | way0Age_103; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2805 = _GEN_4853 | way0Age_104; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2806 = _GEN_4854 | way0Age_105; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2807 = _GEN_4855 | way0Age_106; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2808 = _GEN_4856 | way0Age_107; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2809 = _GEN_4857 | way0Age_108; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2810 = _GEN_4858 | way0Age_109; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2811 = _GEN_4859 | way0Age_110; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2812 = _GEN_4860 | way0Age_111; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2813 = _GEN_4861 | way0Age_112; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2814 = _GEN_4862 | way0Age_113; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2815 = _GEN_4863 | way0Age_114; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2816 = _GEN_4864 | way0Age_115; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2817 = _GEN_4865 | way0Age_116; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2818 = _GEN_4866 | way0Age_117; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2819 = _GEN_4867 | way0Age_118; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2820 = _GEN_4868 | way0Age_119; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2821 = _GEN_4869 | way0Age_120; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2822 = _GEN_4870 | way0Age_121; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2823 = _GEN_4871 | way0Age_122; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2824 = _GEN_4872 | way0Age_123; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2825 = _GEN_4873 | way0Age_124; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2826 = _GEN_4874 | way0Age_125; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2827 = _GEN_4875 | way0Age_126; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2828 = _GEN_4876 | way0Age_127; // @[DCache.scala 201:{23,23} 36:26]
  wire  _GEN_2957 = _GEN_4749 | way1V_0; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_2958 = _GEN_4750 | way1V_1; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_2959 = _GEN_4751 | way1V_2; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_2960 = _GEN_4752 | way1V_3; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_2961 = _GEN_4753 | way1V_4; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_2962 = _GEN_4754 | way1V_5; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_2963 = _GEN_4755 | way1V_6; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_2964 = _GEN_4756 | way1V_7; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_2965 = _GEN_4757 | way1V_8; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_2966 = _GEN_4758 | way1V_9; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_2967 = _GEN_4759 | way1V_10; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_2968 = _GEN_4760 | way1V_11; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_2969 = _GEN_4761 | way1V_12; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_2970 = _GEN_4762 | way1V_13; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_2971 = _GEN_4763 | way1V_14; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_2972 = _GEN_4764 | way1V_15; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_2973 = _GEN_4765 | way1V_16; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_2974 = _GEN_4766 | way1V_17; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_2975 = _GEN_4767 | way1V_18; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_2976 = _GEN_4768 | way1V_19; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_2977 = _GEN_4769 | way1V_20; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_2978 = _GEN_4770 | way1V_21; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_2979 = _GEN_4771 | way1V_22; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_2980 = _GEN_4772 | way1V_23; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_2981 = _GEN_4773 | way1V_24; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_2982 = _GEN_4774 | way1V_25; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_2983 = _GEN_4775 | way1V_26; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_2984 = _GEN_4776 | way1V_27; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_2985 = _GEN_4777 | way1V_28; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_2986 = _GEN_4778 | way1V_29; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_2987 = _GEN_4779 | way1V_30; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_2988 = _GEN_4780 | way1V_31; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_2989 = _GEN_4781 | way1V_32; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_2990 = _GEN_4782 | way1V_33; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_2991 = _GEN_4783 | way1V_34; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_2992 = _GEN_4784 | way1V_35; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_2993 = _GEN_4785 | way1V_36; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_2994 = _GEN_4786 | way1V_37; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_2995 = _GEN_4787 | way1V_38; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_2996 = _GEN_4788 | way1V_39; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_2997 = _GEN_4789 | way1V_40; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_2998 = _GEN_4790 | way1V_41; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_2999 = _GEN_4791 | way1V_42; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_3000 = _GEN_4792 | way1V_43; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_3001 = _GEN_4793 | way1V_44; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_3002 = _GEN_4794 | way1V_45; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_3003 = _GEN_4795 | way1V_46; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_3004 = _GEN_4796 | way1V_47; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_3005 = _GEN_4797 | way1V_48; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_3006 = _GEN_4798 | way1V_49; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_3007 = _GEN_4799 | way1V_50; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_3008 = _GEN_4800 | way1V_51; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_3009 = _GEN_4801 | way1V_52; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_3010 = _GEN_4802 | way1V_53; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_3011 = _GEN_4803 | way1V_54; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_3012 = _GEN_4804 | way1V_55; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_3013 = _GEN_4805 | way1V_56; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_3014 = _GEN_4806 | way1V_57; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_3015 = _GEN_4807 | way1V_58; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_3016 = _GEN_4808 | way1V_59; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_3017 = _GEN_4809 | way1V_60; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_3018 = _GEN_4810 | way1V_61; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_3019 = _GEN_4811 | way1V_62; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_3020 = _GEN_4812 | way1V_63; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_3021 = _GEN_4813 | way1V_64; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_3022 = _GEN_4814 | way1V_65; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_3023 = _GEN_4815 | way1V_66; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_3024 = _GEN_4816 | way1V_67; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_3025 = _GEN_4817 | way1V_68; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_3026 = _GEN_4818 | way1V_69; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_3027 = _GEN_4819 | way1V_70; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_3028 = _GEN_4820 | way1V_71; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_3029 = _GEN_4821 | way1V_72; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_3030 = _GEN_4822 | way1V_73; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_3031 = _GEN_4823 | way1V_74; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_3032 = _GEN_4824 | way1V_75; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_3033 = _GEN_4825 | way1V_76; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_3034 = _GEN_4826 | way1V_77; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_3035 = _GEN_4827 | way1V_78; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_3036 = _GEN_4828 | way1V_79; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_3037 = _GEN_4829 | way1V_80; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_3038 = _GEN_4830 | way1V_81; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_3039 = _GEN_4831 | way1V_82; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_3040 = _GEN_4832 | way1V_83; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_3041 = _GEN_4833 | way1V_84; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_3042 = _GEN_4834 | way1V_85; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_3043 = _GEN_4835 | way1V_86; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_3044 = _GEN_4836 | way1V_87; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_3045 = _GEN_4837 | way1V_88; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_3046 = _GEN_4838 | way1V_89; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_3047 = _GEN_4839 | way1V_90; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_3048 = _GEN_4840 | way1V_91; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_3049 = _GEN_4841 | way1V_92; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_3050 = _GEN_4842 | way1V_93; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_3051 = _GEN_4843 | way1V_94; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_3052 = _GEN_4844 | way1V_95; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_3053 = _GEN_4845 | way1V_96; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_3054 = _GEN_4846 | way1V_97; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_3055 = _GEN_4847 | way1V_98; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_3056 = _GEN_4848 | way1V_99; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_3057 = _GEN_4849 | way1V_100; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_3058 = _GEN_4850 | way1V_101; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_3059 = _GEN_4851 | way1V_102; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_3060 = _GEN_4852 | way1V_103; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_3061 = _GEN_4853 | way1V_104; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_3062 = _GEN_4854 | way1V_105; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_3063 = _GEN_4855 | way1V_106; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_3064 = _GEN_4856 | way1V_107; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_3065 = _GEN_4857 | way1V_108; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_3066 = _GEN_4858 | way1V_109; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_3067 = _GEN_4859 | way1V_110; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_3068 = _GEN_4860 | way1V_111; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_3069 = _GEN_4861 | way1V_112; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_3070 = _GEN_4862 | way1V_113; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_3071 = _GEN_4863 | way1V_114; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_3072 = _GEN_4864 | way1V_115; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_3073 = _GEN_4865 | way1V_116; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_3074 = _GEN_4866 | way1V_117; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_3075 = _GEN_4867 | way1V_118; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_3076 = _GEN_4868 | way1V_119; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_3077 = _GEN_4869 | way1V_120; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_3078 = _GEN_4870 | way1V_121; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_3079 = _GEN_4871 | way1V_122; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_3080 = _GEN_4872 | way1V_123; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_3081 = _GEN_4873 | way1V_124; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_3082 = _GEN_4874 | way1V_125; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_3083 = _GEN_4875 | way1V_126; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_3084 = _GEN_4876 | way1V_127; // @[DCache.scala 204:{21,21} 39:26]
  wire  _GEN_3341 = _GEN_4749 | way1Age_0; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3342 = _GEN_4750 | way1Age_1; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3343 = _GEN_4751 | way1Age_2; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3344 = _GEN_4752 | way1Age_3; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3345 = _GEN_4753 | way1Age_4; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3346 = _GEN_4754 | way1Age_5; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3347 = _GEN_4755 | way1Age_6; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3348 = _GEN_4756 | way1Age_7; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3349 = _GEN_4757 | way1Age_8; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3350 = _GEN_4758 | way1Age_9; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3351 = _GEN_4759 | way1Age_10; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3352 = _GEN_4760 | way1Age_11; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3353 = _GEN_4761 | way1Age_12; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3354 = _GEN_4762 | way1Age_13; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3355 = _GEN_4763 | way1Age_14; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3356 = _GEN_4764 | way1Age_15; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3357 = _GEN_4765 | way1Age_16; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3358 = _GEN_4766 | way1Age_17; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3359 = _GEN_4767 | way1Age_18; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3360 = _GEN_4768 | way1Age_19; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3361 = _GEN_4769 | way1Age_20; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3362 = _GEN_4770 | way1Age_21; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3363 = _GEN_4771 | way1Age_22; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3364 = _GEN_4772 | way1Age_23; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3365 = _GEN_4773 | way1Age_24; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3366 = _GEN_4774 | way1Age_25; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3367 = _GEN_4775 | way1Age_26; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3368 = _GEN_4776 | way1Age_27; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3369 = _GEN_4777 | way1Age_28; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3370 = _GEN_4778 | way1Age_29; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3371 = _GEN_4779 | way1Age_30; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3372 = _GEN_4780 | way1Age_31; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3373 = _GEN_4781 | way1Age_32; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3374 = _GEN_4782 | way1Age_33; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3375 = _GEN_4783 | way1Age_34; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3376 = _GEN_4784 | way1Age_35; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3377 = _GEN_4785 | way1Age_36; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3378 = _GEN_4786 | way1Age_37; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3379 = _GEN_4787 | way1Age_38; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3380 = _GEN_4788 | way1Age_39; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3381 = _GEN_4789 | way1Age_40; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3382 = _GEN_4790 | way1Age_41; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3383 = _GEN_4791 | way1Age_42; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3384 = _GEN_4792 | way1Age_43; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3385 = _GEN_4793 | way1Age_44; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3386 = _GEN_4794 | way1Age_45; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3387 = _GEN_4795 | way1Age_46; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3388 = _GEN_4796 | way1Age_47; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3389 = _GEN_4797 | way1Age_48; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3390 = _GEN_4798 | way1Age_49; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3391 = _GEN_4799 | way1Age_50; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3392 = _GEN_4800 | way1Age_51; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3393 = _GEN_4801 | way1Age_52; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3394 = _GEN_4802 | way1Age_53; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3395 = _GEN_4803 | way1Age_54; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3396 = _GEN_4804 | way1Age_55; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3397 = _GEN_4805 | way1Age_56; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3398 = _GEN_4806 | way1Age_57; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3399 = _GEN_4807 | way1Age_58; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3400 = _GEN_4808 | way1Age_59; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3401 = _GEN_4809 | way1Age_60; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3402 = _GEN_4810 | way1Age_61; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3403 = _GEN_4811 | way1Age_62; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3404 = _GEN_4812 | way1Age_63; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3405 = _GEN_4813 | way1Age_64; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3406 = _GEN_4814 | way1Age_65; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3407 = _GEN_4815 | way1Age_66; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3408 = _GEN_4816 | way1Age_67; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3409 = _GEN_4817 | way1Age_68; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3410 = _GEN_4818 | way1Age_69; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3411 = _GEN_4819 | way1Age_70; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3412 = _GEN_4820 | way1Age_71; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3413 = _GEN_4821 | way1Age_72; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3414 = _GEN_4822 | way1Age_73; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3415 = _GEN_4823 | way1Age_74; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3416 = _GEN_4824 | way1Age_75; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3417 = _GEN_4825 | way1Age_76; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3418 = _GEN_4826 | way1Age_77; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3419 = _GEN_4827 | way1Age_78; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3420 = _GEN_4828 | way1Age_79; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3421 = _GEN_4829 | way1Age_80; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3422 = _GEN_4830 | way1Age_81; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3423 = _GEN_4831 | way1Age_82; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3424 = _GEN_4832 | way1Age_83; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3425 = _GEN_4833 | way1Age_84; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3426 = _GEN_4834 | way1Age_85; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3427 = _GEN_4835 | way1Age_86; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3428 = _GEN_4836 | way1Age_87; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3429 = _GEN_4837 | way1Age_88; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3430 = _GEN_4838 | way1Age_89; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3431 = _GEN_4839 | way1Age_90; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3432 = _GEN_4840 | way1Age_91; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3433 = _GEN_4841 | way1Age_92; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3434 = _GEN_4842 | way1Age_93; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3435 = _GEN_4843 | way1Age_94; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3436 = _GEN_4844 | way1Age_95; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3437 = _GEN_4845 | way1Age_96; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3438 = _GEN_4846 | way1Age_97; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3439 = _GEN_4847 | way1Age_98; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3440 = _GEN_4848 | way1Age_99; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3441 = _GEN_4849 | way1Age_100; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3442 = _GEN_4850 | way1Age_101; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3443 = _GEN_4851 | way1Age_102; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3444 = _GEN_4852 | way1Age_103; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3445 = _GEN_4853 | way1Age_104; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3446 = _GEN_4854 | way1Age_105; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3447 = _GEN_4855 | way1Age_106; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3448 = _GEN_4856 | way1Age_107; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3449 = _GEN_4857 | way1Age_108; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3450 = _GEN_4858 | way1Age_109; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3451 = _GEN_4859 | way1Age_110; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3452 = _GEN_4860 | way1Age_111; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3453 = _GEN_4861 | way1Age_112; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3454 = _GEN_4862 | way1Age_113; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3455 = _GEN_4863 | way1Age_114; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3456 = _GEN_4864 | way1Age_115; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3457 = _GEN_4865 | way1Age_116; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3458 = _GEN_4866 | way1Age_117; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3459 = _GEN_4867 | way1Age_118; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3460 = _GEN_4868 | way1Age_119; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3461 = _GEN_4869 | way1Age_120; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3462 = _GEN_4870 | way1Age_121; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3463 = _GEN_4871 | way1Age_122; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3464 = _GEN_4872 | way1Age_123; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3465 = _GEN_4873 | way1Age_124; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3466 = _GEN_4874 | way1Age_125; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3467 = _GEN_4875 | way1Age_126; // @[DCache.scala 207:{23,23} 42:26]
  wire  _GEN_3468 = _GEN_4876 | way1Age_127; // @[DCache.scala 207:{23,23} 42:26]
  reg  hitEn; // @[DCache.scala 210:22]
  wire [127:0] _rData_T = sDoneEn ? io_out_data_read : 128'h0; // @[DCache.scala 213:20]
  wire [127:0] rData = hitEn ? cacheRData : _rData_T; // @[DCache.scala 212:18]
  wire [63:0] rDataHL = reqOff[3] ? rData[127:64] : rData[63:0]; // @[DCache.scala 214:20]
  wire [7:0] _io_dmem_data_read_T_10 = 3'h1 == reqOff[2:0] ? rDataHL[15:8] : rDataHL[7:0]; // @[Mux.scala 81:58]
  wire [7:0] _io_dmem_data_read_T_12 = 3'h2 == reqOff[2:0] ? rDataHL[23:16] : _io_dmem_data_read_T_10; // @[Mux.scala 81:58]
  wire [7:0] _io_dmem_data_read_T_14 = 3'h3 == reqOff[2:0] ? rDataHL[31:24] : _io_dmem_data_read_T_12; // @[Mux.scala 81:58]
  wire [7:0] _io_dmem_data_read_T_16 = 3'h4 == reqOff[2:0] ? rDataHL[39:32] : _io_dmem_data_read_T_14; // @[Mux.scala 81:58]
  wire [7:0] _io_dmem_data_read_T_18 = 3'h5 == reqOff[2:0] ? rDataHL[47:40] : _io_dmem_data_read_T_16; // @[Mux.scala 81:58]
  wire [7:0] _io_dmem_data_read_T_20 = 3'h6 == reqOff[2:0] ? rDataHL[55:48] : _io_dmem_data_read_T_18; // @[Mux.scala 81:58]
  wire [7:0] _io_dmem_data_read_T_22 = 3'h7 == reqOff[2:0] ? rDataHL[63:56] : _io_dmem_data_read_T_20; // @[Mux.scala 81:58]
  wire [15:0] _io_dmem_data_read_T_29 = 2'h1 == reqOff[2:1] ? rDataHL[31:16] : rDataHL[15:0]; // @[Mux.scala 81:58]
  wire [15:0] _io_dmem_data_read_T_31 = 2'h2 == reqOff[2:1] ? rDataHL[47:32] : _io_dmem_data_read_T_29; // @[Mux.scala 81:58]
  wire [15:0] _io_dmem_data_read_T_33 = 2'h3 == reqOff[2:1] ? rDataHL[63:48] : _io_dmem_data_read_T_31; // @[Mux.scala 81:58]
  wire [31:0] _io_dmem_data_read_T_38 = reqOff[2] ? rDataHL[63:32] : rDataHL[31:0]; // @[Mux.scala 81:58]
  wire [15:0] _io_dmem_data_read_T_40 = 2'h1 == io_dmem_data_size ? _io_dmem_data_read_T_33 : {{8'd0},
    _io_dmem_data_read_T_22}; // @[Mux.scala 81:58]
  wire [31:0] _io_dmem_data_read_T_42 = 2'h2 == io_dmem_data_size ? _io_dmem_data_read_T_38 : {{16'd0},
    _io_dmem_data_read_T_40}; // @[Mux.scala 81:58]
  wire [31:0] _io_out_data_addr_T_1 = {_GEN_140,reqIndex,4'h0}; // @[Cat.scala 31:58]
  wire [31:0] _io_out_data_addr_T_2 = {_GEN_396,reqIndex,4'h0}; // @[Cat.scala 31:58]
  wire [31:0] _io_out_data_addr_T_3 = _cacheDirtyEn_T ? _io_out_data_addr_T_1 : _io_out_data_addr_T_2; // @[DCache.scala 246:26]
  wire [31:0] _io_out_data_addr_T_5 = {io_dmem_data_addr[31:4],4'h0}; // @[Cat.scala 31:58]
  S011HD1P_X32Y2D128_BW req ( // @[DCache.scala 253:19]
    .Q(req_Q),
    .CLK(req_CLK),
    .CEN(req_CEN),
    .WEN(req_WEN),
    .BWEN(req_BWEN),
    .A(req_A),
    .D(req_D)
  );
  assign io_dmem_data_ready = io_dmem_data_req ? sDoneEn : hitEn | sDoneEn; // @[DCache.scala 216:23]
  assign io_dmem_data_read = 2'h3 == io_dmem_data_size ? rDataHL : {{32'd0}, _io_dmem_data_read_T_42}; // @[Mux.scala 81:58]
  assign io_out_data_valid = sWriteEn | sReadEn; // @[DCache.scala 242:24]
  assign io_out_data_req = state == 3'h3; // @[DCache.scala 138:24]
  assign io_out_data_addr = sWriteEn ? _io_out_data_addr_T_3 : _io_out_data_addr_T_5; // @[DCache.scala 245:24]
  assign io_out_data_strb = sWriteEn ? 8'hff : 8'h0; // @[DCache.scala 249:24]
  assign io_out_data_write = sWriteEn ? cacheRData : 128'h0; // @[DCache.scala 250:24]
  assign req_CLK = clock; // @[DCache.scala 254:14]
  assign req_CEN = 1'h1; // @[DCache.scala 255:14]
  assign req_WEN = sCacheWEn | sReadEn & io_out_data_ready; // @[DCache.scala 175:28]
  assign req_BWEN = _valid_WEn_T ? 128'hffffffffffffffffffffffffffffffff : _valid_BWEn_T_1; // @[DCache.scala 178:21]
  assign req_A = _cacheDirtyEn_T ? _cacheIndex_T_1 : _cacheIndex_T_2; // @[DCache.scala 133:22]
  assign req_D = _valid_WEn_T ? io_out_data_read : _valid_WData_T_1; // @[DCache.scala 176:21]
  always @(posedge clock) begin
    if (reset) begin // @[DCache.scala 33:26]
      way0V_0 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_0 <= _GEN_2445;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_1 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_1 <= _GEN_2446;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_2 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_2 <= _GEN_2447;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_3 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_3 <= _GEN_2448;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_4 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_4 <= _GEN_2449;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_5 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_5 <= _GEN_2450;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_6 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_6 <= _GEN_2451;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_7 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_7 <= _GEN_2452;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_8 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_8 <= _GEN_2453;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_9 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_9 <= _GEN_2454;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_10 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_10 <= _GEN_2455;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_11 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_11 <= _GEN_2456;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_12 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_12 <= _GEN_2457;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_13 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_13 <= _GEN_2458;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_14 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_14 <= _GEN_2459;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_15 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_15 <= _GEN_2460;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_16 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_16 <= _GEN_2461;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_17 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_17 <= _GEN_2462;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_18 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_18 <= _GEN_2463;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_19 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_19 <= _GEN_2464;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_20 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_20 <= _GEN_2465;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_21 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_21 <= _GEN_2466;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_22 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_22 <= _GEN_2467;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_23 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_23 <= _GEN_2468;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_24 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_24 <= _GEN_2469;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_25 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_25 <= _GEN_2470;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_26 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_26 <= _GEN_2471;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_27 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_27 <= _GEN_2472;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_28 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_28 <= _GEN_2473;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_29 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_29 <= _GEN_2474;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_30 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_30 <= _GEN_2475;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_31 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_31 <= _GEN_2476;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_32 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_32 <= _GEN_2477;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_33 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_33 <= _GEN_2478;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_34 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_34 <= _GEN_2479;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_35 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_35 <= _GEN_2480;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_36 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_36 <= _GEN_2481;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_37 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_37 <= _GEN_2482;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_38 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_38 <= _GEN_2483;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_39 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_39 <= _GEN_2484;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_40 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_40 <= _GEN_2485;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_41 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_41 <= _GEN_2486;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_42 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_42 <= _GEN_2487;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_43 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_43 <= _GEN_2488;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_44 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_44 <= _GEN_2489;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_45 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_45 <= _GEN_2490;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_46 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_46 <= _GEN_2491;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_47 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_47 <= _GEN_2492;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_48 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_48 <= _GEN_2493;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_49 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_49 <= _GEN_2494;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_50 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_50 <= _GEN_2495;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_51 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_51 <= _GEN_2496;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_52 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_52 <= _GEN_2497;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_53 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_53 <= _GEN_2498;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_54 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_54 <= _GEN_2499;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_55 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_55 <= _GEN_2500;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_56 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_56 <= _GEN_2501;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_57 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_57 <= _GEN_2502;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_58 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_58 <= _GEN_2503;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_59 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_59 <= _GEN_2504;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_60 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_60 <= _GEN_2505;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_61 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_61 <= _GEN_2506;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_62 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_62 <= _GEN_2507;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_63 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_63 <= _GEN_2508;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_64 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_64 <= _GEN_2509;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_65 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_65 <= _GEN_2510;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_66 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_66 <= _GEN_2511;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_67 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_67 <= _GEN_2512;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_68 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_68 <= _GEN_2513;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_69 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_69 <= _GEN_2514;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_70 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_70 <= _GEN_2515;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_71 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_71 <= _GEN_2516;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_72 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_72 <= _GEN_2517;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_73 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_73 <= _GEN_2518;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_74 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_74 <= _GEN_2519;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_75 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_75 <= _GEN_2520;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_76 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_76 <= _GEN_2521;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_77 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_77 <= _GEN_2522;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_78 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_78 <= _GEN_2523;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_79 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_79 <= _GEN_2524;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_80 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_80 <= _GEN_2525;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_81 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_81 <= _GEN_2526;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_82 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_82 <= _GEN_2527;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_83 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_83 <= _GEN_2528;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_84 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_84 <= _GEN_2529;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_85 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_85 <= _GEN_2530;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_86 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_86 <= _GEN_2531;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_87 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_87 <= _GEN_2532;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_88 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_88 <= _GEN_2533;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_89 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_89 <= _GEN_2534;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_90 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_90 <= _GEN_2535;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_91 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_91 <= _GEN_2536;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_92 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_92 <= _GEN_2537;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_93 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_93 <= _GEN_2538;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_94 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_94 <= _GEN_2539;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_95 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_95 <= _GEN_2540;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_96 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_96 <= _GEN_2541;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_97 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_97 <= _GEN_2542;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_98 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_98 <= _GEN_2543;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_99 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_99 <= _GEN_2544;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_100 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_100 <= _GEN_2545;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_101 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_101 <= _GEN_2546;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_102 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_102 <= _GEN_2547;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_103 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_103 <= _GEN_2548;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_104 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_104 <= _GEN_2549;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_105 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_105 <= _GEN_2550;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_106 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_106 <= _GEN_2551;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_107 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_107 <= _GEN_2552;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_108 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_108 <= _GEN_2553;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_109 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_109 <= _GEN_2554;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_110 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_110 <= _GEN_2555;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_111 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_111 <= _GEN_2556;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_112 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_112 <= _GEN_2557;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_113 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_113 <= _GEN_2558;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_114 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_114 <= _GEN_2559;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_115 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_115 <= _GEN_2560;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_116 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_116 <= _GEN_2561;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_117 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_117 <= _GEN_2562;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_118 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_118 <= _GEN_2563;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_119 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_119 <= _GEN_2564;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_120 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_120 <= _GEN_2565;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_121 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_121 <= _GEN_2566;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_122 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_122 <= _GEN_2567;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_123 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_123 <= _GEN_2568;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_124 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_124 <= _GEN_2569;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_125 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_125 <= _GEN_2570;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_126 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_126 <= _GEN_2571;
    end
    if (reset) begin // @[DCache.scala 33:26]
      way0V_127 <= 1'h0; // @[DCache.scala 33:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0V_127 <= _GEN_2572;
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_0 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h0 == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_0 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_1 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h1 == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_1 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_2 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h2 == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_2 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_3 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h3 == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_3 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_4 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h4 == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_4 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_5 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h5 == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_5 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_6 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h6 == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_6 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_7 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h7 == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_7 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_8 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h8 == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_8 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_9 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h9 == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_9 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_10 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'ha == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_10 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_11 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'hb == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_11 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_12 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'hc == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_12 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_13 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'hd == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_13 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_14 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'he == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_14 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_15 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'hf == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_15 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_16 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h10 == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_16 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_17 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h11 == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_17 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_18 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h12 == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_18 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_19 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h13 == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_19 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_20 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h14 == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_20 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_21 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h15 == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_21 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_22 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h16 == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_22 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_23 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h17 == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_23 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_24 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h18 == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_24 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_25 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h19 == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_25 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_26 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h1a == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_26 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_27 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h1b == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_27 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_28 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h1c == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_28 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_29 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h1d == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_29 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_30 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h1e == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_30 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_31 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h1f == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_31 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_32 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h20 == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_32 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_33 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h21 == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_33 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_34 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h22 == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_34 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_35 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h23 == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_35 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_36 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h24 == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_36 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_37 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h25 == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_37 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_38 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h26 == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_38 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_39 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h27 == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_39 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_40 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h28 == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_40 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_41 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h29 == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_41 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_42 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h2a == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_42 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_43 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h2b == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_43 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_44 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h2c == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_44 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_45 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h2d == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_45 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_46 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h2e == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_46 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_47 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h2f == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_47 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_48 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h30 == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_48 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_49 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h31 == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_49 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_50 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h32 == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_50 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_51 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h33 == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_51 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_52 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h34 == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_52 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_53 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h35 == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_53 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_54 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h36 == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_54 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_55 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h37 == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_55 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_56 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h38 == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_56 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_57 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h39 == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_57 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_58 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h3a == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_58 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_59 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h3b == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_59 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_60 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h3c == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_60 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_61 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h3d == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_61 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_62 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h3e == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_62 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_63 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h3f == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_63 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_64 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h40 == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_64 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_65 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h41 == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_65 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_66 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h42 == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_66 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_67 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h43 == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_67 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_68 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h44 == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_68 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_69 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h45 == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_69 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_70 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h46 == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_70 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_71 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h47 == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_71 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_72 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h48 == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_72 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_73 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h49 == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_73 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_74 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h4a == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_74 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_75 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h4b == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_75 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_76 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h4c == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_76 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_77 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h4d == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_77 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_78 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h4e == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_78 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_79 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h4f == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_79 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_80 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h50 == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_80 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_81 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h51 == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_81 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_82 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h52 == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_82 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_83 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h53 == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_83 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_84 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h54 == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_84 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_85 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h55 == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_85 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_86 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h56 == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_86 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_87 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h57 == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_87 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_88 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h58 == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_88 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_89 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h59 == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_89 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_90 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h5a == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_90 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_91 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h5b == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_91 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_92 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h5c == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_92 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_93 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h5d == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_93 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_94 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h5e == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_94 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_95 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h5f == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_95 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_96 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h60 == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_96 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_97 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h61 == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_97 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_98 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h62 == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_98 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_99 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h63 == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_99 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_100 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h64 == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_100 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_101 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h65 == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_101 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_102 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h66 == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_102 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_103 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h67 == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_103 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_104 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h68 == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_104 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_105 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h69 == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_105 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_106 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h6a == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_106 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_107 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h6b == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_107 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_108 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h6c == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_108 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_109 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h6d == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_109 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_110 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h6e == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_110 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_111 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h6f == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_111 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_112 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h70 == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_112 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_113 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h71 == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_113 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_114 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h72 == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_114 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_115 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h73 == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_115 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_116 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h74 == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_116 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_117 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h75 == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_117 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_118 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h76 == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_118 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_119 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h77 == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_119 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_120 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h78 == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_120 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_121 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h79 == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_121 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_122 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h7a == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_122 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_123 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h7b == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_123 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_124 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h7c == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_124 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_125 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h7d == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_125 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_126 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h7e == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_126 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 34:26]
      way0Tag_127 <= 21'h0; // @[DCache.scala 34:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h7f == reqIndex) begin // @[DCache.scala 200:23]
        way0Tag_127 <= reqTag; // @[DCache.scala 200:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_0 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_0 <= _GEN_2701;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h0 == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_0 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_1 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_1 <= _GEN_2702;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h1 == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_1 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_2 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_2 <= _GEN_2703;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h2 == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_2 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_3 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_3 <= _GEN_2704;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h3 == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_3 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_4 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_4 <= _GEN_2705;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h4 == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_4 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_5 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_5 <= _GEN_2706;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h5 == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_5 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_6 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_6 <= _GEN_2707;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h6 == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_6 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_7 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_7 <= _GEN_2708;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h7 == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_7 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_8 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_8 <= _GEN_2709;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h8 == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_8 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_9 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_9 <= _GEN_2710;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h9 == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_9 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_10 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_10 <= _GEN_2711;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'ha == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_10 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_11 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_11 <= _GEN_2712;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'hb == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_11 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_12 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_12 <= _GEN_2713;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'hc == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_12 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_13 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_13 <= _GEN_2714;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'hd == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_13 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_14 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_14 <= _GEN_2715;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'he == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_14 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_15 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_15 <= _GEN_2716;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'hf == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_15 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_16 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_16 <= _GEN_2717;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h10 == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_16 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_17 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_17 <= _GEN_2718;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h11 == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_17 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_18 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_18 <= _GEN_2719;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h12 == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_18 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_19 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_19 <= _GEN_2720;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h13 == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_19 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_20 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_20 <= _GEN_2721;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h14 == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_20 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_21 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_21 <= _GEN_2722;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h15 == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_21 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_22 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_22 <= _GEN_2723;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h16 == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_22 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_23 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_23 <= _GEN_2724;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h17 == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_23 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_24 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_24 <= _GEN_2725;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h18 == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_24 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_25 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_25 <= _GEN_2726;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h19 == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_25 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_26 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_26 <= _GEN_2727;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h1a == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_26 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_27 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_27 <= _GEN_2728;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h1b == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_27 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_28 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_28 <= _GEN_2729;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h1c == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_28 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_29 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_29 <= _GEN_2730;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h1d == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_29 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_30 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_30 <= _GEN_2731;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h1e == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_30 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_31 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_31 <= _GEN_2732;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h1f == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_31 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_32 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_32 <= _GEN_2733;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h20 == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_32 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_33 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_33 <= _GEN_2734;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h21 == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_33 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_34 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_34 <= _GEN_2735;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h22 == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_34 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_35 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_35 <= _GEN_2736;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h23 == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_35 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_36 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_36 <= _GEN_2737;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h24 == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_36 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_37 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_37 <= _GEN_2738;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h25 == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_37 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_38 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_38 <= _GEN_2739;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h26 == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_38 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_39 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_39 <= _GEN_2740;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h27 == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_39 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_40 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_40 <= _GEN_2741;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h28 == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_40 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_41 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_41 <= _GEN_2742;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h29 == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_41 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_42 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_42 <= _GEN_2743;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h2a == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_42 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_43 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_43 <= _GEN_2744;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h2b == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_43 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_44 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_44 <= _GEN_2745;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h2c == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_44 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_45 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_45 <= _GEN_2746;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h2d == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_45 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_46 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_46 <= _GEN_2747;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h2e == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_46 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_47 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_47 <= _GEN_2748;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h2f == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_47 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_48 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_48 <= _GEN_2749;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h30 == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_48 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_49 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_49 <= _GEN_2750;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h31 == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_49 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_50 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_50 <= _GEN_2751;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h32 == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_50 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_51 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_51 <= _GEN_2752;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h33 == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_51 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_52 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_52 <= _GEN_2753;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h34 == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_52 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_53 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_53 <= _GEN_2754;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h35 == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_53 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_54 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_54 <= _GEN_2755;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h36 == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_54 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_55 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_55 <= _GEN_2756;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h37 == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_55 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_56 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_56 <= _GEN_2757;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h38 == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_56 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_57 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_57 <= _GEN_2758;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h39 == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_57 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_58 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_58 <= _GEN_2759;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h3a == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_58 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_59 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_59 <= _GEN_2760;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h3b == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_59 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_60 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_60 <= _GEN_2761;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h3c == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_60 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_61 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_61 <= _GEN_2762;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h3d == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_61 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_62 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_62 <= _GEN_2763;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h3e == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_62 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_63 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_63 <= _GEN_2764;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h3f == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_63 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_64 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_64 <= _GEN_2765;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h40 == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_64 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_65 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_65 <= _GEN_2766;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h41 == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_65 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_66 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_66 <= _GEN_2767;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h42 == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_66 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_67 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_67 <= _GEN_2768;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h43 == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_67 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_68 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_68 <= _GEN_2769;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h44 == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_68 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_69 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_69 <= _GEN_2770;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h45 == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_69 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_70 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_70 <= _GEN_2771;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h46 == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_70 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_71 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_71 <= _GEN_2772;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h47 == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_71 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_72 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_72 <= _GEN_2773;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h48 == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_72 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_73 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_73 <= _GEN_2774;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h49 == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_73 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_74 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_74 <= _GEN_2775;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h4a == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_74 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_75 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_75 <= _GEN_2776;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h4b == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_75 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_76 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_76 <= _GEN_2777;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h4c == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_76 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_77 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_77 <= _GEN_2778;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h4d == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_77 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_78 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_78 <= _GEN_2779;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h4e == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_78 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_79 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_79 <= _GEN_2780;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h4f == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_79 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_80 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_80 <= _GEN_2781;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h50 == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_80 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_81 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_81 <= _GEN_2782;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h51 == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_81 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_82 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_82 <= _GEN_2783;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h52 == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_82 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_83 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_83 <= _GEN_2784;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h53 == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_83 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_84 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_84 <= _GEN_2785;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h54 == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_84 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_85 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_85 <= _GEN_2786;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h55 == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_85 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_86 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_86 <= _GEN_2787;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h56 == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_86 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_87 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_87 <= _GEN_2788;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h57 == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_87 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_88 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_88 <= _GEN_2789;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h58 == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_88 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_89 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_89 <= _GEN_2790;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h59 == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_89 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_90 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_90 <= _GEN_2791;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h5a == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_90 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_91 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_91 <= _GEN_2792;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h5b == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_91 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_92 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_92 <= _GEN_2793;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h5c == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_92 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_93 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_93 <= _GEN_2794;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h5d == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_93 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_94 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_94 <= _GEN_2795;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h5e == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_94 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_95 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_95 <= _GEN_2796;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h5f == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_95 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_96 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_96 <= _GEN_2797;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h60 == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_96 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_97 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_97 <= _GEN_2798;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h61 == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_97 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_98 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_98 <= _GEN_2799;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h62 == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_98 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_99 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_99 <= _GEN_2800;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h63 == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_99 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_100 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_100 <= _GEN_2801;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h64 == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_100 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_101 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_101 <= _GEN_2802;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h65 == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_101 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_102 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_102 <= _GEN_2803;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h66 == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_102 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_103 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_103 <= _GEN_2804;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h67 == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_103 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_104 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_104 <= _GEN_2805;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h68 == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_104 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_105 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_105 <= _GEN_2806;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h69 == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_105 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_106 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_106 <= _GEN_2807;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h6a == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_106 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_107 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_107 <= _GEN_2808;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h6b == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_107 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_108 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_108 <= _GEN_2809;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h6c == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_108 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_109 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_109 <= _GEN_2810;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h6d == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_109 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_110 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_110 <= _GEN_2811;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h6e == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_110 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_111 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_111 <= _GEN_2812;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h6f == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_111 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_112 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_112 <= _GEN_2813;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h70 == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_112 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_113 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_113 <= _GEN_2814;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h71 == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_113 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_114 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_114 <= _GEN_2815;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h72 == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_114 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_115 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_115 <= _GEN_2816;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h73 == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_115 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_116 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_116 <= _GEN_2817;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h74 == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_116 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_117 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_117 <= _GEN_2818;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h75 == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_117 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_118 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_118 <= _GEN_2819;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h76 == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_118 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_119 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_119 <= _GEN_2820;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h77 == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_119 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_120 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_120 <= _GEN_2821;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h78 == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_120 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_121 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_121 <= _GEN_2822;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h79 == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_121 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_122 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_122 <= _GEN_2823;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h7a == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_122 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_123 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_123 <= _GEN_2824;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h7b == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_123 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_124 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_124 <= _GEN_2825;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h7c == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_124 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_125 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_125 <= _GEN_2826;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h7d == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_125 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_126 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_126 <= _GEN_2827;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h7e == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_126 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 36:26]
      way0Age_127 <= 1'h0; // @[DCache.scala 36:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      way0Age_127 <= _GEN_2828;
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      if (7'h7f == reqIndex) begin // @[DCache.scala 206:23]
        way0Age_127 <= 1'h0; // @[DCache.scala 206:23]
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_0 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_0 <= _GEN_1037;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_0 <= _GEN_1165;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_1 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_1 <= _GEN_1038;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_1 <= _GEN_1166;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_2 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_2 <= _GEN_1039;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_2 <= _GEN_1167;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_3 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_3 <= _GEN_1040;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_3 <= _GEN_1168;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_4 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_4 <= _GEN_1041;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_4 <= _GEN_1169;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_5 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_5 <= _GEN_1042;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_5 <= _GEN_1170;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_6 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_6 <= _GEN_1043;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_6 <= _GEN_1171;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_7 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_7 <= _GEN_1044;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_7 <= _GEN_1172;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_8 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_8 <= _GEN_1045;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_8 <= _GEN_1173;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_9 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_9 <= _GEN_1046;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_9 <= _GEN_1174;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_10 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_10 <= _GEN_1047;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_10 <= _GEN_1175;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_11 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_11 <= _GEN_1048;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_11 <= _GEN_1176;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_12 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_12 <= _GEN_1049;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_12 <= _GEN_1177;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_13 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_13 <= _GEN_1050;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_13 <= _GEN_1178;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_14 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_14 <= _GEN_1051;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_14 <= _GEN_1179;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_15 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_15 <= _GEN_1052;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_15 <= _GEN_1180;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_16 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_16 <= _GEN_1053;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_16 <= _GEN_1181;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_17 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_17 <= _GEN_1054;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_17 <= _GEN_1182;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_18 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_18 <= _GEN_1055;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_18 <= _GEN_1183;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_19 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_19 <= _GEN_1056;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_19 <= _GEN_1184;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_20 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_20 <= _GEN_1057;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_20 <= _GEN_1185;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_21 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_21 <= _GEN_1058;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_21 <= _GEN_1186;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_22 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_22 <= _GEN_1059;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_22 <= _GEN_1187;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_23 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_23 <= _GEN_1060;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_23 <= _GEN_1188;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_24 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_24 <= _GEN_1061;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_24 <= _GEN_1189;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_25 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_25 <= _GEN_1062;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_25 <= _GEN_1190;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_26 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_26 <= _GEN_1063;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_26 <= _GEN_1191;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_27 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_27 <= _GEN_1064;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_27 <= _GEN_1192;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_28 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_28 <= _GEN_1065;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_28 <= _GEN_1193;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_29 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_29 <= _GEN_1066;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_29 <= _GEN_1194;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_30 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_30 <= _GEN_1067;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_30 <= _GEN_1195;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_31 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_31 <= _GEN_1068;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_31 <= _GEN_1196;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_32 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_32 <= _GEN_1069;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_32 <= _GEN_1197;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_33 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_33 <= _GEN_1070;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_33 <= _GEN_1198;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_34 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_34 <= _GEN_1071;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_34 <= _GEN_1199;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_35 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_35 <= _GEN_1072;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_35 <= _GEN_1200;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_36 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_36 <= _GEN_1073;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_36 <= _GEN_1201;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_37 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_37 <= _GEN_1074;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_37 <= _GEN_1202;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_38 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_38 <= _GEN_1075;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_38 <= _GEN_1203;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_39 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_39 <= _GEN_1076;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_39 <= _GEN_1204;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_40 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_40 <= _GEN_1077;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_40 <= _GEN_1205;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_41 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_41 <= _GEN_1078;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_41 <= _GEN_1206;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_42 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_42 <= _GEN_1079;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_42 <= _GEN_1207;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_43 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_43 <= _GEN_1080;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_43 <= _GEN_1208;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_44 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_44 <= _GEN_1081;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_44 <= _GEN_1209;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_45 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_45 <= _GEN_1082;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_45 <= _GEN_1210;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_46 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_46 <= _GEN_1083;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_46 <= _GEN_1211;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_47 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_47 <= _GEN_1084;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_47 <= _GEN_1212;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_48 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_48 <= _GEN_1085;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_48 <= _GEN_1213;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_49 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_49 <= _GEN_1086;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_49 <= _GEN_1214;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_50 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_50 <= _GEN_1087;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_50 <= _GEN_1215;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_51 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_51 <= _GEN_1088;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_51 <= _GEN_1216;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_52 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_52 <= _GEN_1089;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_52 <= _GEN_1217;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_53 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_53 <= _GEN_1090;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_53 <= _GEN_1218;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_54 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_54 <= _GEN_1091;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_54 <= _GEN_1219;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_55 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_55 <= _GEN_1092;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_55 <= _GEN_1220;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_56 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_56 <= _GEN_1093;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_56 <= _GEN_1221;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_57 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_57 <= _GEN_1094;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_57 <= _GEN_1222;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_58 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_58 <= _GEN_1095;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_58 <= _GEN_1223;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_59 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_59 <= _GEN_1096;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_59 <= _GEN_1224;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_60 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_60 <= _GEN_1097;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_60 <= _GEN_1225;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_61 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_61 <= _GEN_1098;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_61 <= _GEN_1226;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_62 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_62 <= _GEN_1099;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_62 <= _GEN_1227;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_63 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_63 <= _GEN_1100;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_63 <= _GEN_1228;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_64 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_64 <= _GEN_1101;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_64 <= _GEN_1229;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_65 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_65 <= _GEN_1102;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_65 <= _GEN_1230;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_66 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_66 <= _GEN_1103;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_66 <= _GEN_1231;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_67 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_67 <= _GEN_1104;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_67 <= _GEN_1232;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_68 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_68 <= _GEN_1105;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_68 <= _GEN_1233;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_69 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_69 <= _GEN_1106;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_69 <= _GEN_1234;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_70 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_70 <= _GEN_1107;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_70 <= _GEN_1235;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_71 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_71 <= _GEN_1108;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_71 <= _GEN_1236;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_72 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_72 <= _GEN_1109;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_72 <= _GEN_1237;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_73 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_73 <= _GEN_1110;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_73 <= _GEN_1238;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_74 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_74 <= _GEN_1111;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_74 <= _GEN_1239;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_75 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_75 <= _GEN_1112;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_75 <= _GEN_1240;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_76 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_76 <= _GEN_1113;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_76 <= _GEN_1241;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_77 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_77 <= _GEN_1114;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_77 <= _GEN_1242;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_78 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_78 <= _GEN_1115;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_78 <= _GEN_1243;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_79 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_79 <= _GEN_1116;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_79 <= _GEN_1244;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_80 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_80 <= _GEN_1117;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_80 <= _GEN_1245;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_81 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_81 <= _GEN_1118;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_81 <= _GEN_1246;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_82 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_82 <= _GEN_1119;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_82 <= _GEN_1247;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_83 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_83 <= _GEN_1120;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_83 <= _GEN_1248;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_84 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_84 <= _GEN_1121;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_84 <= _GEN_1249;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_85 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_85 <= _GEN_1122;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_85 <= _GEN_1250;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_86 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_86 <= _GEN_1123;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_86 <= _GEN_1251;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_87 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_87 <= _GEN_1124;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_87 <= _GEN_1252;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_88 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_88 <= _GEN_1125;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_88 <= _GEN_1253;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_89 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_89 <= _GEN_1126;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_89 <= _GEN_1254;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_90 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_90 <= _GEN_1127;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_90 <= _GEN_1255;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_91 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_91 <= _GEN_1128;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_91 <= _GEN_1256;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_92 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_92 <= _GEN_1129;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_92 <= _GEN_1257;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_93 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_93 <= _GEN_1130;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_93 <= _GEN_1258;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_94 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_94 <= _GEN_1131;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_94 <= _GEN_1259;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_95 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_95 <= _GEN_1132;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_95 <= _GEN_1260;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_96 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_96 <= _GEN_1133;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_96 <= _GEN_1261;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_97 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_97 <= _GEN_1134;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_97 <= _GEN_1262;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_98 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_98 <= _GEN_1135;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_98 <= _GEN_1263;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_99 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_99 <= _GEN_1136;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_99 <= _GEN_1264;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_100 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_100 <= _GEN_1137;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_100 <= _GEN_1265;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_101 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_101 <= _GEN_1138;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_101 <= _GEN_1266;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_102 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_102 <= _GEN_1139;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_102 <= _GEN_1267;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_103 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_103 <= _GEN_1140;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_103 <= _GEN_1268;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_104 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_104 <= _GEN_1141;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_104 <= _GEN_1269;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_105 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_105 <= _GEN_1142;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_105 <= _GEN_1270;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_106 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_106 <= _GEN_1143;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_106 <= _GEN_1271;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_107 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_107 <= _GEN_1144;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_107 <= _GEN_1272;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_108 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_108 <= _GEN_1145;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_108 <= _GEN_1273;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_109 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_109 <= _GEN_1146;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_109 <= _GEN_1274;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_110 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_110 <= _GEN_1147;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_110 <= _GEN_1275;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_111 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_111 <= _GEN_1148;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_111 <= _GEN_1276;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_112 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_112 <= _GEN_1149;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_112 <= _GEN_1277;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_113 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_113 <= _GEN_1150;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_113 <= _GEN_1278;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_114 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_114 <= _GEN_1151;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_114 <= _GEN_1279;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_115 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_115 <= _GEN_1152;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_115 <= _GEN_1280;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_116 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_116 <= _GEN_1153;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_116 <= _GEN_1281;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_117 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_117 <= _GEN_1154;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_117 <= _GEN_1282;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_118 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_118 <= _GEN_1155;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_118 <= _GEN_1283;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_119 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_119 <= _GEN_1156;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_119 <= _GEN_1284;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_120 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_120 <= _GEN_1157;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_120 <= _GEN_1285;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_121 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_121 <= _GEN_1158;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_121 <= _GEN_1286;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_122 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_122 <= _GEN_1159;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_122 <= _GEN_1287;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_123 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_123 <= _GEN_1160;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_123 <= _GEN_1288;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_124 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_124 <= _GEN_1161;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_124 <= _GEN_1289;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_125 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_125 <= _GEN_1162;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_125 <= _GEN_1290;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_126 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_126 <= _GEN_1163;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_126 <= _GEN_1291;
      end
    end
    if (reset) begin // @[DCache.scala 37:26]
      way0Dirty_127 <= 1'h0; // @[DCache.scala 37:26]
    end else if (ageWay0En | way0Hit) begin // @[DCache.scala 182:30]
      if (sCacheWEn & io_dmem_data_req) begin // @[DCache.scala 183:36]
        way0Dirty_127 <= _GEN_1164;
      end else if (sWriteEn & io_out_data_ready) begin // @[DCache.scala 185:45]
        way0Dirty_127 <= _GEN_1292;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_0 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_0 <= _GEN_2957;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_1 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_1 <= _GEN_2958;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_2 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_2 <= _GEN_2959;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_3 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_3 <= _GEN_2960;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_4 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_4 <= _GEN_2961;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_5 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_5 <= _GEN_2962;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_6 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_6 <= _GEN_2963;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_7 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_7 <= _GEN_2964;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_8 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_8 <= _GEN_2965;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_9 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_9 <= _GEN_2966;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_10 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_10 <= _GEN_2967;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_11 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_11 <= _GEN_2968;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_12 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_12 <= _GEN_2969;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_13 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_13 <= _GEN_2970;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_14 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_14 <= _GEN_2971;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_15 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_15 <= _GEN_2972;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_16 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_16 <= _GEN_2973;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_17 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_17 <= _GEN_2974;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_18 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_18 <= _GEN_2975;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_19 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_19 <= _GEN_2976;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_20 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_20 <= _GEN_2977;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_21 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_21 <= _GEN_2978;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_22 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_22 <= _GEN_2979;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_23 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_23 <= _GEN_2980;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_24 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_24 <= _GEN_2981;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_25 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_25 <= _GEN_2982;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_26 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_26 <= _GEN_2983;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_27 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_27 <= _GEN_2984;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_28 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_28 <= _GEN_2985;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_29 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_29 <= _GEN_2986;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_30 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_30 <= _GEN_2987;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_31 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_31 <= _GEN_2988;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_32 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_32 <= _GEN_2989;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_33 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_33 <= _GEN_2990;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_34 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_34 <= _GEN_2991;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_35 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_35 <= _GEN_2992;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_36 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_36 <= _GEN_2993;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_37 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_37 <= _GEN_2994;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_38 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_38 <= _GEN_2995;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_39 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_39 <= _GEN_2996;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_40 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_40 <= _GEN_2997;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_41 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_41 <= _GEN_2998;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_42 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_42 <= _GEN_2999;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_43 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_43 <= _GEN_3000;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_44 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_44 <= _GEN_3001;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_45 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_45 <= _GEN_3002;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_46 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_46 <= _GEN_3003;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_47 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_47 <= _GEN_3004;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_48 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_48 <= _GEN_3005;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_49 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_49 <= _GEN_3006;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_50 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_50 <= _GEN_3007;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_51 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_51 <= _GEN_3008;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_52 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_52 <= _GEN_3009;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_53 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_53 <= _GEN_3010;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_54 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_54 <= _GEN_3011;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_55 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_55 <= _GEN_3012;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_56 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_56 <= _GEN_3013;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_57 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_57 <= _GEN_3014;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_58 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_58 <= _GEN_3015;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_59 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_59 <= _GEN_3016;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_60 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_60 <= _GEN_3017;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_61 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_61 <= _GEN_3018;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_62 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_62 <= _GEN_3019;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_63 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_63 <= _GEN_3020;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_64 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_64 <= _GEN_3021;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_65 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_65 <= _GEN_3022;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_66 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_66 <= _GEN_3023;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_67 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_67 <= _GEN_3024;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_68 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_68 <= _GEN_3025;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_69 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_69 <= _GEN_3026;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_70 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_70 <= _GEN_3027;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_71 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_71 <= _GEN_3028;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_72 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_72 <= _GEN_3029;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_73 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_73 <= _GEN_3030;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_74 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_74 <= _GEN_3031;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_75 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_75 <= _GEN_3032;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_76 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_76 <= _GEN_3033;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_77 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_77 <= _GEN_3034;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_78 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_78 <= _GEN_3035;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_79 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_79 <= _GEN_3036;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_80 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_80 <= _GEN_3037;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_81 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_81 <= _GEN_3038;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_82 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_82 <= _GEN_3039;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_83 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_83 <= _GEN_3040;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_84 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_84 <= _GEN_3041;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_85 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_85 <= _GEN_3042;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_86 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_86 <= _GEN_3043;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_87 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_87 <= _GEN_3044;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_88 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_88 <= _GEN_3045;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_89 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_89 <= _GEN_3046;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_90 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_90 <= _GEN_3047;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_91 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_91 <= _GEN_3048;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_92 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_92 <= _GEN_3049;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_93 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_93 <= _GEN_3050;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_94 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_94 <= _GEN_3051;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_95 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_95 <= _GEN_3052;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_96 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_96 <= _GEN_3053;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_97 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_97 <= _GEN_3054;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_98 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_98 <= _GEN_3055;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_99 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_99 <= _GEN_3056;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_100 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_100 <= _GEN_3057;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_101 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_101 <= _GEN_3058;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_102 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_102 <= _GEN_3059;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_103 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_103 <= _GEN_3060;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_104 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_104 <= _GEN_3061;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_105 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_105 <= _GEN_3062;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_106 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_106 <= _GEN_3063;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_107 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_107 <= _GEN_3064;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_108 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_108 <= _GEN_3065;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_109 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_109 <= _GEN_3066;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_110 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_110 <= _GEN_3067;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_111 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_111 <= _GEN_3068;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_112 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_112 <= _GEN_3069;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_113 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_113 <= _GEN_3070;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_114 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_114 <= _GEN_3071;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_115 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_115 <= _GEN_3072;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_116 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_116 <= _GEN_3073;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_117 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_117 <= _GEN_3074;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_118 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_118 <= _GEN_3075;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_119 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_119 <= _GEN_3076;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_120 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_120 <= _GEN_3077;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_121 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_121 <= _GEN_3078;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_122 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_122 <= _GEN_3079;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_123 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_123 <= _GEN_3080;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_124 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_124 <= _GEN_3081;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_125 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_125 <= _GEN_3082;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_126 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_126 <= _GEN_3083;
      end
    end
    if (reset) begin // @[DCache.scala 39:26]
      way1V_127 <= 1'h0; // @[DCache.scala 39:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        way1V_127 <= _GEN_3084;
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_0 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h0 == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_0 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_1 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h1 == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_1 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_2 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h2 == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_2 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_3 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h3 == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_3 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_4 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h4 == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_4 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_5 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h5 == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_5 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_6 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h6 == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_6 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_7 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h7 == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_7 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_8 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h8 == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_8 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_9 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h9 == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_9 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_10 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'ha == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_10 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_11 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'hb == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_11 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_12 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'hc == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_12 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_13 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'hd == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_13 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_14 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'he == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_14 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_15 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'hf == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_15 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_16 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h10 == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_16 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_17 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h11 == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_17 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_18 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h12 == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_18 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_19 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h13 == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_19 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_20 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h14 == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_20 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_21 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h15 == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_21 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_22 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h16 == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_22 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_23 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h17 == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_23 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_24 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h18 == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_24 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_25 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h19 == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_25 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_26 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h1a == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_26 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_27 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h1b == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_27 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_28 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h1c == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_28 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_29 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h1d == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_29 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_30 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h1e == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_30 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_31 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h1f == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_31 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_32 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h20 == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_32 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_33 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h21 == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_33 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_34 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h22 == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_34 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_35 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h23 == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_35 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_36 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h24 == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_36 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_37 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h25 == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_37 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_38 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h26 == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_38 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_39 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h27 == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_39 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_40 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h28 == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_40 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_41 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h29 == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_41 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_42 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h2a == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_42 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_43 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h2b == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_43 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_44 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h2c == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_44 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_45 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h2d == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_45 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_46 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h2e == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_46 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_47 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h2f == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_47 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_48 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h30 == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_48 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_49 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h31 == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_49 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_50 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h32 == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_50 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_51 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h33 == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_51 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_52 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h34 == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_52 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_53 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h35 == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_53 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_54 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h36 == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_54 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_55 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h37 == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_55 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_56 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h38 == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_56 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_57 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h39 == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_57 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_58 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h3a == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_58 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_59 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h3b == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_59 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_60 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h3c == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_60 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_61 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h3d == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_61 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_62 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h3e == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_62 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_63 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h3f == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_63 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_64 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h40 == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_64 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_65 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h41 == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_65 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_66 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h42 == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_66 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_67 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h43 == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_67 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_68 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h44 == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_68 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_69 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h45 == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_69 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_70 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h46 == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_70 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_71 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h47 == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_71 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_72 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h48 == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_72 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_73 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h49 == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_73 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_74 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h4a == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_74 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_75 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h4b == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_75 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_76 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h4c == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_76 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_77 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h4d == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_77 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_78 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h4e == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_78 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_79 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h4f == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_79 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_80 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h50 == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_80 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_81 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h51 == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_81 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_82 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h52 == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_82 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_83 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h53 == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_83 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_84 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h54 == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_84 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_85 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h55 == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_85 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_86 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h56 == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_86 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_87 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h57 == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_87 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_88 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h58 == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_88 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_89 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h59 == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_89 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_90 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h5a == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_90 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_91 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h5b == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_91 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_92 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h5c == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_92 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_93 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h5d == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_93 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_94 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h5e == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_94 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_95 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h5f == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_95 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_96 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h60 == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_96 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_97 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h61 == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_97 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_98 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h62 == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_98 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_99 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h63 == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_99 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_100 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h64 == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_100 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_101 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h65 == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_101 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_102 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h66 == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_102 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_103 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h67 == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_103 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_104 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h68 == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_104 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_105 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h69 == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_105 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_106 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h6a == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_106 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_107 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h6b == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_107 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_108 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h6c == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_108 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_109 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h6d == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_109 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_110 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h6e == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_110 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_111 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h6f == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_111 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_112 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h70 == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_112 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_113 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h71 == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_113 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_114 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h72 == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_114 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_115 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h73 == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_115 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_116 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h74 == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_116 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_117 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h75 == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_117 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_118 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h76 == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_118 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_119 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h77 == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_119 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_120 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h78 == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_120 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_121 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h79 == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_121 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_122 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h7a == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_122 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_123 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h7b == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_123 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_124 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h7c == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_124 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_125 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h7d == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_125 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_126 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h7e == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_126 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 40:26]
      way1Tag_127 <= 21'h0; // @[DCache.scala 40:26]
    end else if (!(ageWay0En & sDoneEn)) begin // @[DCache.scala 198:30]
      if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
        if (7'h7f == reqIndex) begin // @[DCache.scala 205:23]
          way1Tag_127 <= reqTag; // @[DCache.scala 205:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_0 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h0 == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_0 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_0 <= _GEN_3341;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_1 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h1 == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_1 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_1 <= _GEN_3342;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_2 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h2 == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_2 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_2 <= _GEN_3343;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_3 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h3 == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_3 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_3 <= _GEN_3344;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_4 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h4 == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_4 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_4 <= _GEN_3345;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_5 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h5 == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_5 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_5 <= _GEN_3346;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_6 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h6 == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_6 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_6 <= _GEN_3347;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_7 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h7 == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_7 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_7 <= _GEN_3348;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_8 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h8 == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_8 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_8 <= _GEN_3349;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_9 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h9 == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_9 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_9 <= _GEN_3350;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_10 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'ha == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_10 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_10 <= _GEN_3351;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_11 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'hb == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_11 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_11 <= _GEN_3352;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_12 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'hc == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_12 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_12 <= _GEN_3353;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_13 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'hd == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_13 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_13 <= _GEN_3354;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_14 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'he == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_14 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_14 <= _GEN_3355;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_15 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'hf == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_15 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_15 <= _GEN_3356;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_16 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h10 == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_16 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_16 <= _GEN_3357;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_17 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h11 == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_17 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_17 <= _GEN_3358;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_18 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h12 == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_18 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_18 <= _GEN_3359;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_19 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h13 == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_19 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_19 <= _GEN_3360;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_20 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h14 == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_20 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_20 <= _GEN_3361;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_21 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h15 == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_21 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_21 <= _GEN_3362;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_22 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h16 == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_22 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_22 <= _GEN_3363;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_23 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h17 == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_23 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_23 <= _GEN_3364;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_24 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h18 == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_24 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_24 <= _GEN_3365;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_25 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h19 == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_25 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_25 <= _GEN_3366;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_26 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h1a == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_26 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_26 <= _GEN_3367;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_27 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h1b == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_27 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_27 <= _GEN_3368;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_28 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h1c == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_28 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_28 <= _GEN_3369;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_29 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h1d == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_29 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_29 <= _GEN_3370;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_30 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h1e == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_30 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_30 <= _GEN_3371;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_31 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h1f == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_31 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_31 <= _GEN_3372;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_32 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h20 == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_32 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_32 <= _GEN_3373;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_33 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h21 == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_33 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_33 <= _GEN_3374;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_34 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h22 == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_34 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_34 <= _GEN_3375;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_35 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h23 == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_35 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_35 <= _GEN_3376;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_36 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h24 == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_36 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_36 <= _GEN_3377;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_37 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h25 == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_37 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_37 <= _GEN_3378;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_38 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h26 == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_38 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_38 <= _GEN_3379;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_39 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h27 == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_39 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_39 <= _GEN_3380;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_40 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h28 == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_40 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_40 <= _GEN_3381;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_41 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h29 == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_41 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_41 <= _GEN_3382;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_42 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h2a == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_42 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_42 <= _GEN_3383;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_43 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h2b == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_43 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_43 <= _GEN_3384;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_44 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h2c == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_44 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_44 <= _GEN_3385;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_45 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h2d == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_45 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_45 <= _GEN_3386;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_46 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h2e == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_46 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_46 <= _GEN_3387;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_47 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h2f == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_47 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_47 <= _GEN_3388;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_48 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h30 == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_48 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_48 <= _GEN_3389;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_49 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h31 == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_49 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_49 <= _GEN_3390;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_50 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h32 == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_50 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_50 <= _GEN_3391;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_51 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h33 == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_51 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_51 <= _GEN_3392;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_52 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h34 == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_52 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_52 <= _GEN_3393;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_53 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h35 == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_53 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_53 <= _GEN_3394;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_54 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h36 == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_54 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_54 <= _GEN_3395;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_55 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h37 == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_55 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_55 <= _GEN_3396;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_56 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h38 == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_56 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_56 <= _GEN_3397;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_57 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h39 == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_57 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_57 <= _GEN_3398;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_58 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h3a == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_58 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_58 <= _GEN_3399;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_59 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h3b == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_59 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_59 <= _GEN_3400;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_60 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h3c == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_60 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_60 <= _GEN_3401;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_61 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h3d == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_61 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_61 <= _GEN_3402;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_62 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h3e == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_62 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_62 <= _GEN_3403;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_63 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h3f == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_63 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_63 <= _GEN_3404;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_64 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h40 == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_64 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_64 <= _GEN_3405;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_65 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h41 == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_65 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_65 <= _GEN_3406;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_66 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h42 == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_66 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_66 <= _GEN_3407;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_67 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h43 == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_67 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_67 <= _GEN_3408;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_68 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h44 == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_68 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_68 <= _GEN_3409;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_69 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h45 == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_69 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_69 <= _GEN_3410;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_70 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h46 == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_70 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_70 <= _GEN_3411;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_71 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h47 == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_71 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_71 <= _GEN_3412;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_72 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h48 == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_72 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_72 <= _GEN_3413;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_73 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h49 == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_73 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_73 <= _GEN_3414;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_74 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h4a == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_74 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_74 <= _GEN_3415;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_75 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h4b == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_75 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_75 <= _GEN_3416;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_76 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h4c == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_76 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_76 <= _GEN_3417;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_77 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h4d == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_77 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_77 <= _GEN_3418;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_78 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h4e == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_78 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_78 <= _GEN_3419;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_79 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h4f == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_79 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_79 <= _GEN_3420;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_80 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h50 == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_80 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_80 <= _GEN_3421;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_81 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h51 == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_81 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_81 <= _GEN_3422;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_82 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h52 == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_82 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_82 <= _GEN_3423;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_83 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h53 == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_83 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_83 <= _GEN_3424;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_84 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h54 == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_84 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_84 <= _GEN_3425;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_85 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h55 == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_85 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_85 <= _GEN_3426;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_86 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h56 == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_86 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_86 <= _GEN_3427;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_87 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h57 == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_87 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_87 <= _GEN_3428;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_88 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h58 == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_88 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_88 <= _GEN_3429;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_89 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h59 == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_89 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_89 <= _GEN_3430;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_90 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h5a == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_90 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_90 <= _GEN_3431;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_91 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h5b == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_91 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_91 <= _GEN_3432;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_92 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h5c == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_92 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_92 <= _GEN_3433;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_93 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h5d == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_93 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_93 <= _GEN_3434;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_94 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h5e == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_94 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_94 <= _GEN_3435;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_95 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h5f == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_95 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_95 <= _GEN_3436;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_96 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h60 == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_96 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_96 <= _GEN_3437;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_97 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h61 == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_97 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_97 <= _GEN_3438;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_98 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h62 == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_98 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_98 <= _GEN_3439;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_99 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h63 == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_99 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_99 <= _GEN_3440;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_100 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h64 == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_100 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_100 <= _GEN_3441;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_101 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h65 == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_101 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_101 <= _GEN_3442;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_102 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h66 == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_102 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_102 <= _GEN_3443;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_103 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h67 == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_103 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_103 <= _GEN_3444;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_104 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h68 == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_104 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_104 <= _GEN_3445;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_105 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h69 == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_105 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_105 <= _GEN_3446;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_106 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h6a == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_106 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_106 <= _GEN_3447;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_107 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h6b == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_107 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_107 <= _GEN_3448;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_108 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h6c == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_108 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_108 <= _GEN_3449;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_109 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h6d == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_109 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_109 <= _GEN_3450;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_110 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h6e == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_110 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_110 <= _GEN_3451;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_111 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h6f == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_111 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_111 <= _GEN_3452;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_112 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h70 == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_112 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_112 <= _GEN_3453;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_113 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h71 == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_113 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_113 <= _GEN_3454;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_114 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h72 == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_114 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_114 <= _GEN_3455;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_115 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h73 == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_115 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_115 <= _GEN_3456;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_116 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h74 == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_116 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_116 <= _GEN_3457;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_117 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h75 == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_117 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_117 <= _GEN_3458;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_118 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h76 == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_118 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_118 <= _GEN_3459;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_119 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h77 == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_119 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_119 <= _GEN_3460;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_120 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h78 == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_120 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_120 <= _GEN_3461;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_121 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h79 == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_121 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_121 <= _GEN_3462;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_122 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h7a == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_122 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_122 <= _GEN_3463;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_123 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h7b == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_123 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_123 <= _GEN_3464;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_124 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h7c == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_124 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_124 <= _GEN_3465;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_125 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h7d == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_125 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_125 <= _GEN_3466;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_126 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h7e == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_126 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_126 <= _GEN_3467;
    end
    if (reset) begin // @[DCache.scala 42:26]
      way1Age_127 <= 1'h0; // @[DCache.scala 42:26]
    end else if (ageWay0En & sDoneEn) begin // @[DCache.scala 198:30]
      if (7'h7f == reqIndex) begin // @[DCache.scala 202:23]
        way1Age_127 <= 1'h0; // @[DCache.scala 202:23]
      end
    end else if (ageWay1En & sDoneEn) begin // @[DCache.scala 203:37]
      way1Age_127 <= _GEN_3468;
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_0 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_0 <= _GEN_1549;
        end else begin
          way1Dirty_0 <= _GEN_1805;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_1 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_1 <= _GEN_1550;
        end else begin
          way1Dirty_1 <= _GEN_1806;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_2 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_2 <= _GEN_1551;
        end else begin
          way1Dirty_2 <= _GEN_1807;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_3 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_3 <= _GEN_1552;
        end else begin
          way1Dirty_3 <= _GEN_1808;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_4 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_4 <= _GEN_1553;
        end else begin
          way1Dirty_4 <= _GEN_1809;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_5 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_5 <= _GEN_1554;
        end else begin
          way1Dirty_5 <= _GEN_1810;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_6 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_6 <= _GEN_1555;
        end else begin
          way1Dirty_6 <= _GEN_1811;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_7 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_7 <= _GEN_1556;
        end else begin
          way1Dirty_7 <= _GEN_1812;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_8 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_8 <= _GEN_1557;
        end else begin
          way1Dirty_8 <= _GEN_1813;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_9 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_9 <= _GEN_1558;
        end else begin
          way1Dirty_9 <= _GEN_1814;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_10 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_10 <= _GEN_1559;
        end else begin
          way1Dirty_10 <= _GEN_1815;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_11 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_11 <= _GEN_1560;
        end else begin
          way1Dirty_11 <= _GEN_1816;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_12 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_12 <= _GEN_1561;
        end else begin
          way1Dirty_12 <= _GEN_1817;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_13 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_13 <= _GEN_1562;
        end else begin
          way1Dirty_13 <= _GEN_1818;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_14 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_14 <= _GEN_1563;
        end else begin
          way1Dirty_14 <= _GEN_1819;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_15 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_15 <= _GEN_1564;
        end else begin
          way1Dirty_15 <= _GEN_1820;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_16 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_16 <= _GEN_1565;
        end else begin
          way1Dirty_16 <= _GEN_1821;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_17 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_17 <= _GEN_1566;
        end else begin
          way1Dirty_17 <= _GEN_1822;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_18 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_18 <= _GEN_1567;
        end else begin
          way1Dirty_18 <= _GEN_1823;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_19 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_19 <= _GEN_1568;
        end else begin
          way1Dirty_19 <= _GEN_1824;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_20 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_20 <= _GEN_1569;
        end else begin
          way1Dirty_20 <= _GEN_1825;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_21 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_21 <= _GEN_1570;
        end else begin
          way1Dirty_21 <= _GEN_1826;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_22 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_22 <= _GEN_1571;
        end else begin
          way1Dirty_22 <= _GEN_1827;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_23 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_23 <= _GEN_1572;
        end else begin
          way1Dirty_23 <= _GEN_1828;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_24 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_24 <= _GEN_1573;
        end else begin
          way1Dirty_24 <= _GEN_1829;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_25 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_25 <= _GEN_1574;
        end else begin
          way1Dirty_25 <= _GEN_1830;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_26 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_26 <= _GEN_1575;
        end else begin
          way1Dirty_26 <= _GEN_1831;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_27 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_27 <= _GEN_1576;
        end else begin
          way1Dirty_27 <= _GEN_1832;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_28 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_28 <= _GEN_1577;
        end else begin
          way1Dirty_28 <= _GEN_1833;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_29 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_29 <= _GEN_1578;
        end else begin
          way1Dirty_29 <= _GEN_1834;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_30 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_30 <= _GEN_1579;
        end else begin
          way1Dirty_30 <= _GEN_1835;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_31 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_31 <= _GEN_1580;
        end else begin
          way1Dirty_31 <= _GEN_1836;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_32 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_32 <= _GEN_1581;
        end else begin
          way1Dirty_32 <= _GEN_1837;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_33 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_33 <= _GEN_1582;
        end else begin
          way1Dirty_33 <= _GEN_1838;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_34 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_34 <= _GEN_1583;
        end else begin
          way1Dirty_34 <= _GEN_1839;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_35 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_35 <= _GEN_1584;
        end else begin
          way1Dirty_35 <= _GEN_1840;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_36 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_36 <= _GEN_1585;
        end else begin
          way1Dirty_36 <= _GEN_1841;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_37 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_37 <= _GEN_1586;
        end else begin
          way1Dirty_37 <= _GEN_1842;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_38 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_38 <= _GEN_1587;
        end else begin
          way1Dirty_38 <= _GEN_1843;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_39 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_39 <= _GEN_1588;
        end else begin
          way1Dirty_39 <= _GEN_1844;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_40 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_40 <= _GEN_1589;
        end else begin
          way1Dirty_40 <= _GEN_1845;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_41 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_41 <= _GEN_1590;
        end else begin
          way1Dirty_41 <= _GEN_1846;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_42 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_42 <= _GEN_1591;
        end else begin
          way1Dirty_42 <= _GEN_1847;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_43 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_43 <= _GEN_1592;
        end else begin
          way1Dirty_43 <= _GEN_1848;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_44 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_44 <= _GEN_1593;
        end else begin
          way1Dirty_44 <= _GEN_1849;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_45 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_45 <= _GEN_1594;
        end else begin
          way1Dirty_45 <= _GEN_1850;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_46 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_46 <= _GEN_1595;
        end else begin
          way1Dirty_46 <= _GEN_1851;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_47 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_47 <= _GEN_1596;
        end else begin
          way1Dirty_47 <= _GEN_1852;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_48 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_48 <= _GEN_1597;
        end else begin
          way1Dirty_48 <= _GEN_1853;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_49 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_49 <= _GEN_1598;
        end else begin
          way1Dirty_49 <= _GEN_1854;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_50 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_50 <= _GEN_1599;
        end else begin
          way1Dirty_50 <= _GEN_1855;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_51 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_51 <= _GEN_1600;
        end else begin
          way1Dirty_51 <= _GEN_1856;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_52 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_52 <= _GEN_1601;
        end else begin
          way1Dirty_52 <= _GEN_1857;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_53 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_53 <= _GEN_1602;
        end else begin
          way1Dirty_53 <= _GEN_1858;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_54 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_54 <= _GEN_1603;
        end else begin
          way1Dirty_54 <= _GEN_1859;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_55 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_55 <= _GEN_1604;
        end else begin
          way1Dirty_55 <= _GEN_1860;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_56 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_56 <= _GEN_1605;
        end else begin
          way1Dirty_56 <= _GEN_1861;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_57 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_57 <= _GEN_1606;
        end else begin
          way1Dirty_57 <= _GEN_1862;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_58 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_58 <= _GEN_1607;
        end else begin
          way1Dirty_58 <= _GEN_1863;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_59 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_59 <= _GEN_1608;
        end else begin
          way1Dirty_59 <= _GEN_1864;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_60 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_60 <= _GEN_1609;
        end else begin
          way1Dirty_60 <= _GEN_1865;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_61 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_61 <= _GEN_1610;
        end else begin
          way1Dirty_61 <= _GEN_1866;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_62 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_62 <= _GEN_1611;
        end else begin
          way1Dirty_62 <= _GEN_1867;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_63 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_63 <= _GEN_1612;
        end else begin
          way1Dirty_63 <= _GEN_1868;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_64 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_64 <= _GEN_1613;
        end else begin
          way1Dirty_64 <= _GEN_1869;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_65 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_65 <= _GEN_1614;
        end else begin
          way1Dirty_65 <= _GEN_1870;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_66 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_66 <= _GEN_1615;
        end else begin
          way1Dirty_66 <= _GEN_1871;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_67 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_67 <= _GEN_1616;
        end else begin
          way1Dirty_67 <= _GEN_1872;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_68 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_68 <= _GEN_1617;
        end else begin
          way1Dirty_68 <= _GEN_1873;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_69 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_69 <= _GEN_1618;
        end else begin
          way1Dirty_69 <= _GEN_1874;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_70 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_70 <= _GEN_1619;
        end else begin
          way1Dirty_70 <= _GEN_1875;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_71 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_71 <= _GEN_1620;
        end else begin
          way1Dirty_71 <= _GEN_1876;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_72 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_72 <= _GEN_1621;
        end else begin
          way1Dirty_72 <= _GEN_1877;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_73 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_73 <= _GEN_1622;
        end else begin
          way1Dirty_73 <= _GEN_1878;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_74 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_74 <= _GEN_1623;
        end else begin
          way1Dirty_74 <= _GEN_1879;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_75 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_75 <= _GEN_1624;
        end else begin
          way1Dirty_75 <= _GEN_1880;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_76 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_76 <= _GEN_1625;
        end else begin
          way1Dirty_76 <= _GEN_1881;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_77 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_77 <= _GEN_1626;
        end else begin
          way1Dirty_77 <= _GEN_1882;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_78 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_78 <= _GEN_1627;
        end else begin
          way1Dirty_78 <= _GEN_1883;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_79 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_79 <= _GEN_1628;
        end else begin
          way1Dirty_79 <= _GEN_1884;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_80 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_80 <= _GEN_1629;
        end else begin
          way1Dirty_80 <= _GEN_1885;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_81 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_81 <= _GEN_1630;
        end else begin
          way1Dirty_81 <= _GEN_1886;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_82 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_82 <= _GEN_1631;
        end else begin
          way1Dirty_82 <= _GEN_1887;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_83 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_83 <= _GEN_1632;
        end else begin
          way1Dirty_83 <= _GEN_1888;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_84 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_84 <= _GEN_1633;
        end else begin
          way1Dirty_84 <= _GEN_1889;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_85 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_85 <= _GEN_1634;
        end else begin
          way1Dirty_85 <= _GEN_1890;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_86 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_86 <= _GEN_1635;
        end else begin
          way1Dirty_86 <= _GEN_1891;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_87 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_87 <= _GEN_1636;
        end else begin
          way1Dirty_87 <= _GEN_1892;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_88 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_88 <= _GEN_1637;
        end else begin
          way1Dirty_88 <= _GEN_1893;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_89 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_89 <= _GEN_1638;
        end else begin
          way1Dirty_89 <= _GEN_1894;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_90 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_90 <= _GEN_1639;
        end else begin
          way1Dirty_90 <= _GEN_1895;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_91 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_91 <= _GEN_1640;
        end else begin
          way1Dirty_91 <= _GEN_1896;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_92 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_92 <= _GEN_1641;
        end else begin
          way1Dirty_92 <= _GEN_1897;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_93 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_93 <= _GEN_1642;
        end else begin
          way1Dirty_93 <= _GEN_1898;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_94 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_94 <= _GEN_1643;
        end else begin
          way1Dirty_94 <= _GEN_1899;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_95 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_95 <= _GEN_1644;
        end else begin
          way1Dirty_95 <= _GEN_1900;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_96 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_96 <= _GEN_1645;
        end else begin
          way1Dirty_96 <= _GEN_1901;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_97 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_97 <= _GEN_1646;
        end else begin
          way1Dirty_97 <= _GEN_1902;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_98 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_98 <= _GEN_1647;
        end else begin
          way1Dirty_98 <= _GEN_1903;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_99 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_99 <= _GEN_1648;
        end else begin
          way1Dirty_99 <= _GEN_1904;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_100 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_100 <= _GEN_1649;
        end else begin
          way1Dirty_100 <= _GEN_1905;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_101 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_101 <= _GEN_1650;
        end else begin
          way1Dirty_101 <= _GEN_1906;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_102 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_102 <= _GEN_1651;
        end else begin
          way1Dirty_102 <= _GEN_1907;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_103 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_103 <= _GEN_1652;
        end else begin
          way1Dirty_103 <= _GEN_1908;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_104 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_104 <= _GEN_1653;
        end else begin
          way1Dirty_104 <= _GEN_1909;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_105 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_105 <= _GEN_1654;
        end else begin
          way1Dirty_105 <= _GEN_1910;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_106 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_106 <= _GEN_1655;
        end else begin
          way1Dirty_106 <= _GEN_1911;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_107 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_107 <= _GEN_1656;
        end else begin
          way1Dirty_107 <= _GEN_1912;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_108 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_108 <= _GEN_1657;
        end else begin
          way1Dirty_108 <= _GEN_1913;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_109 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_109 <= _GEN_1658;
        end else begin
          way1Dirty_109 <= _GEN_1914;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_110 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_110 <= _GEN_1659;
        end else begin
          way1Dirty_110 <= _GEN_1915;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_111 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_111 <= _GEN_1660;
        end else begin
          way1Dirty_111 <= _GEN_1916;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_112 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_112 <= _GEN_1661;
        end else begin
          way1Dirty_112 <= _GEN_1917;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_113 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_113 <= _GEN_1662;
        end else begin
          way1Dirty_113 <= _GEN_1918;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_114 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_114 <= _GEN_1663;
        end else begin
          way1Dirty_114 <= _GEN_1919;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_115 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_115 <= _GEN_1664;
        end else begin
          way1Dirty_115 <= _GEN_1920;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_116 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_116 <= _GEN_1665;
        end else begin
          way1Dirty_116 <= _GEN_1921;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_117 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_117 <= _GEN_1666;
        end else begin
          way1Dirty_117 <= _GEN_1922;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_118 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_118 <= _GEN_1667;
        end else begin
          way1Dirty_118 <= _GEN_1923;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_119 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_119 <= _GEN_1668;
        end else begin
          way1Dirty_119 <= _GEN_1924;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_120 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_120 <= _GEN_1669;
        end else begin
          way1Dirty_120 <= _GEN_1925;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_121 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_121 <= _GEN_1670;
        end else begin
          way1Dirty_121 <= _GEN_1926;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_122 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_122 <= _GEN_1671;
        end else begin
          way1Dirty_122 <= _GEN_1927;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_123 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_123 <= _GEN_1672;
        end else begin
          way1Dirty_123 <= _GEN_1928;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_124 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_124 <= _GEN_1673;
        end else begin
          way1Dirty_124 <= _GEN_1929;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_125 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_125 <= _GEN_1674;
        end else begin
          way1Dirty_125 <= _GEN_1930;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_126 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_126 <= _GEN_1675;
        end else begin
          way1Dirty_126 <= _GEN_1931;
        end
      end
    end
    if (reset) begin // @[DCache.scala 43:26]
      way1Dirty_127 <= 1'h0; // @[DCache.scala 43:26]
    end else if (!(ageWay0En | way0Hit)) begin // @[DCache.scala 182:30]
      if (ageWay1En | way1Hit) begin // @[DCache.scala 188:37]
        if (_T_9) begin // @[DCache.scala 189:36]
          way1Dirty_127 <= _GEN_1676;
        end else begin
          way1Dirty_127 <= _GEN_1932;
        end
      end
    end
    if (reset) begin // @[DCache.scala 46:22]
      state <= 3'h0; // @[DCache.scala 46:22]
    end else if (3'h0 == state) begin // @[DCache.scala 77:17]
      if (io_dmem_data_valid) begin // @[DCache.scala 79:25]
        state <= 3'h1; // @[DCache.scala 80:15]
      end
    end else if (3'h1 == state) begin // @[DCache.scala 77:17]
      if (cacheHitEn) begin // @[DCache.scala 84:27]
        state <= _GEN_1;
      end else begin
        state <= 3'h2; // @[DCache.scala 91:15]
      end
    end else if (3'h2 == state) begin // @[DCache.scala 77:17]
      state <= _GEN_3;
    end else begin
      state <= _GEN_9;
    end
    if (reset) begin // @[DCache.scala 210:22]
      hitEn <= 1'h0; // @[DCache.scala 210:22]
    end else begin
      hitEn <= sHitEn & cacheHitEn; // @[DCache.scala 211:9]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  way0V_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  way0V_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  way0V_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  way0V_3 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  way0V_4 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  way0V_5 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  way0V_6 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  way0V_7 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  way0V_8 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  way0V_9 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  way0V_10 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  way0V_11 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  way0V_12 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  way0V_13 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  way0V_14 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  way0V_15 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  way0V_16 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  way0V_17 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  way0V_18 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  way0V_19 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  way0V_20 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  way0V_21 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  way0V_22 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  way0V_23 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  way0V_24 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  way0V_25 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  way0V_26 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  way0V_27 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  way0V_28 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  way0V_29 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  way0V_30 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  way0V_31 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  way0V_32 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  way0V_33 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  way0V_34 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  way0V_35 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  way0V_36 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  way0V_37 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  way0V_38 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  way0V_39 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  way0V_40 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  way0V_41 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  way0V_42 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  way0V_43 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  way0V_44 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  way0V_45 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  way0V_46 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  way0V_47 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  way0V_48 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  way0V_49 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  way0V_50 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  way0V_51 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  way0V_52 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  way0V_53 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  way0V_54 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  way0V_55 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  way0V_56 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  way0V_57 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  way0V_58 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  way0V_59 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  way0V_60 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  way0V_61 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  way0V_62 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  way0V_63 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  way0V_64 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  way0V_65 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  way0V_66 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  way0V_67 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  way0V_68 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  way0V_69 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  way0V_70 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  way0V_71 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  way0V_72 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  way0V_73 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  way0V_74 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  way0V_75 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  way0V_76 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  way0V_77 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  way0V_78 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  way0V_79 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  way0V_80 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  way0V_81 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  way0V_82 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  way0V_83 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  way0V_84 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  way0V_85 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  way0V_86 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  way0V_87 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  way0V_88 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  way0V_89 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  way0V_90 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  way0V_91 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  way0V_92 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  way0V_93 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  way0V_94 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  way0V_95 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  way0V_96 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  way0V_97 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  way0V_98 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  way0V_99 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  way0V_100 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  way0V_101 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  way0V_102 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  way0V_103 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  way0V_104 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  way0V_105 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  way0V_106 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  way0V_107 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  way0V_108 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  way0V_109 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  way0V_110 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  way0V_111 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  way0V_112 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  way0V_113 = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  way0V_114 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  way0V_115 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  way0V_116 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  way0V_117 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  way0V_118 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  way0V_119 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  way0V_120 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  way0V_121 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  way0V_122 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  way0V_123 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  way0V_124 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  way0V_125 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  way0V_126 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  way0V_127 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  way0Tag_0 = _RAND_128[20:0];
  _RAND_129 = {1{`RANDOM}};
  way0Tag_1 = _RAND_129[20:0];
  _RAND_130 = {1{`RANDOM}};
  way0Tag_2 = _RAND_130[20:0];
  _RAND_131 = {1{`RANDOM}};
  way0Tag_3 = _RAND_131[20:0];
  _RAND_132 = {1{`RANDOM}};
  way0Tag_4 = _RAND_132[20:0];
  _RAND_133 = {1{`RANDOM}};
  way0Tag_5 = _RAND_133[20:0];
  _RAND_134 = {1{`RANDOM}};
  way0Tag_6 = _RAND_134[20:0];
  _RAND_135 = {1{`RANDOM}};
  way0Tag_7 = _RAND_135[20:0];
  _RAND_136 = {1{`RANDOM}};
  way0Tag_8 = _RAND_136[20:0];
  _RAND_137 = {1{`RANDOM}};
  way0Tag_9 = _RAND_137[20:0];
  _RAND_138 = {1{`RANDOM}};
  way0Tag_10 = _RAND_138[20:0];
  _RAND_139 = {1{`RANDOM}};
  way0Tag_11 = _RAND_139[20:0];
  _RAND_140 = {1{`RANDOM}};
  way0Tag_12 = _RAND_140[20:0];
  _RAND_141 = {1{`RANDOM}};
  way0Tag_13 = _RAND_141[20:0];
  _RAND_142 = {1{`RANDOM}};
  way0Tag_14 = _RAND_142[20:0];
  _RAND_143 = {1{`RANDOM}};
  way0Tag_15 = _RAND_143[20:0];
  _RAND_144 = {1{`RANDOM}};
  way0Tag_16 = _RAND_144[20:0];
  _RAND_145 = {1{`RANDOM}};
  way0Tag_17 = _RAND_145[20:0];
  _RAND_146 = {1{`RANDOM}};
  way0Tag_18 = _RAND_146[20:0];
  _RAND_147 = {1{`RANDOM}};
  way0Tag_19 = _RAND_147[20:0];
  _RAND_148 = {1{`RANDOM}};
  way0Tag_20 = _RAND_148[20:0];
  _RAND_149 = {1{`RANDOM}};
  way0Tag_21 = _RAND_149[20:0];
  _RAND_150 = {1{`RANDOM}};
  way0Tag_22 = _RAND_150[20:0];
  _RAND_151 = {1{`RANDOM}};
  way0Tag_23 = _RAND_151[20:0];
  _RAND_152 = {1{`RANDOM}};
  way0Tag_24 = _RAND_152[20:0];
  _RAND_153 = {1{`RANDOM}};
  way0Tag_25 = _RAND_153[20:0];
  _RAND_154 = {1{`RANDOM}};
  way0Tag_26 = _RAND_154[20:0];
  _RAND_155 = {1{`RANDOM}};
  way0Tag_27 = _RAND_155[20:0];
  _RAND_156 = {1{`RANDOM}};
  way0Tag_28 = _RAND_156[20:0];
  _RAND_157 = {1{`RANDOM}};
  way0Tag_29 = _RAND_157[20:0];
  _RAND_158 = {1{`RANDOM}};
  way0Tag_30 = _RAND_158[20:0];
  _RAND_159 = {1{`RANDOM}};
  way0Tag_31 = _RAND_159[20:0];
  _RAND_160 = {1{`RANDOM}};
  way0Tag_32 = _RAND_160[20:0];
  _RAND_161 = {1{`RANDOM}};
  way0Tag_33 = _RAND_161[20:0];
  _RAND_162 = {1{`RANDOM}};
  way0Tag_34 = _RAND_162[20:0];
  _RAND_163 = {1{`RANDOM}};
  way0Tag_35 = _RAND_163[20:0];
  _RAND_164 = {1{`RANDOM}};
  way0Tag_36 = _RAND_164[20:0];
  _RAND_165 = {1{`RANDOM}};
  way0Tag_37 = _RAND_165[20:0];
  _RAND_166 = {1{`RANDOM}};
  way0Tag_38 = _RAND_166[20:0];
  _RAND_167 = {1{`RANDOM}};
  way0Tag_39 = _RAND_167[20:0];
  _RAND_168 = {1{`RANDOM}};
  way0Tag_40 = _RAND_168[20:0];
  _RAND_169 = {1{`RANDOM}};
  way0Tag_41 = _RAND_169[20:0];
  _RAND_170 = {1{`RANDOM}};
  way0Tag_42 = _RAND_170[20:0];
  _RAND_171 = {1{`RANDOM}};
  way0Tag_43 = _RAND_171[20:0];
  _RAND_172 = {1{`RANDOM}};
  way0Tag_44 = _RAND_172[20:0];
  _RAND_173 = {1{`RANDOM}};
  way0Tag_45 = _RAND_173[20:0];
  _RAND_174 = {1{`RANDOM}};
  way0Tag_46 = _RAND_174[20:0];
  _RAND_175 = {1{`RANDOM}};
  way0Tag_47 = _RAND_175[20:0];
  _RAND_176 = {1{`RANDOM}};
  way0Tag_48 = _RAND_176[20:0];
  _RAND_177 = {1{`RANDOM}};
  way0Tag_49 = _RAND_177[20:0];
  _RAND_178 = {1{`RANDOM}};
  way0Tag_50 = _RAND_178[20:0];
  _RAND_179 = {1{`RANDOM}};
  way0Tag_51 = _RAND_179[20:0];
  _RAND_180 = {1{`RANDOM}};
  way0Tag_52 = _RAND_180[20:0];
  _RAND_181 = {1{`RANDOM}};
  way0Tag_53 = _RAND_181[20:0];
  _RAND_182 = {1{`RANDOM}};
  way0Tag_54 = _RAND_182[20:0];
  _RAND_183 = {1{`RANDOM}};
  way0Tag_55 = _RAND_183[20:0];
  _RAND_184 = {1{`RANDOM}};
  way0Tag_56 = _RAND_184[20:0];
  _RAND_185 = {1{`RANDOM}};
  way0Tag_57 = _RAND_185[20:0];
  _RAND_186 = {1{`RANDOM}};
  way0Tag_58 = _RAND_186[20:0];
  _RAND_187 = {1{`RANDOM}};
  way0Tag_59 = _RAND_187[20:0];
  _RAND_188 = {1{`RANDOM}};
  way0Tag_60 = _RAND_188[20:0];
  _RAND_189 = {1{`RANDOM}};
  way0Tag_61 = _RAND_189[20:0];
  _RAND_190 = {1{`RANDOM}};
  way0Tag_62 = _RAND_190[20:0];
  _RAND_191 = {1{`RANDOM}};
  way0Tag_63 = _RAND_191[20:0];
  _RAND_192 = {1{`RANDOM}};
  way0Tag_64 = _RAND_192[20:0];
  _RAND_193 = {1{`RANDOM}};
  way0Tag_65 = _RAND_193[20:0];
  _RAND_194 = {1{`RANDOM}};
  way0Tag_66 = _RAND_194[20:0];
  _RAND_195 = {1{`RANDOM}};
  way0Tag_67 = _RAND_195[20:0];
  _RAND_196 = {1{`RANDOM}};
  way0Tag_68 = _RAND_196[20:0];
  _RAND_197 = {1{`RANDOM}};
  way0Tag_69 = _RAND_197[20:0];
  _RAND_198 = {1{`RANDOM}};
  way0Tag_70 = _RAND_198[20:0];
  _RAND_199 = {1{`RANDOM}};
  way0Tag_71 = _RAND_199[20:0];
  _RAND_200 = {1{`RANDOM}};
  way0Tag_72 = _RAND_200[20:0];
  _RAND_201 = {1{`RANDOM}};
  way0Tag_73 = _RAND_201[20:0];
  _RAND_202 = {1{`RANDOM}};
  way0Tag_74 = _RAND_202[20:0];
  _RAND_203 = {1{`RANDOM}};
  way0Tag_75 = _RAND_203[20:0];
  _RAND_204 = {1{`RANDOM}};
  way0Tag_76 = _RAND_204[20:0];
  _RAND_205 = {1{`RANDOM}};
  way0Tag_77 = _RAND_205[20:0];
  _RAND_206 = {1{`RANDOM}};
  way0Tag_78 = _RAND_206[20:0];
  _RAND_207 = {1{`RANDOM}};
  way0Tag_79 = _RAND_207[20:0];
  _RAND_208 = {1{`RANDOM}};
  way0Tag_80 = _RAND_208[20:0];
  _RAND_209 = {1{`RANDOM}};
  way0Tag_81 = _RAND_209[20:0];
  _RAND_210 = {1{`RANDOM}};
  way0Tag_82 = _RAND_210[20:0];
  _RAND_211 = {1{`RANDOM}};
  way0Tag_83 = _RAND_211[20:0];
  _RAND_212 = {1{`RANDOM}};
  way0Tag_84 = _RAND_212[20:0];
  _RAND_213 = {1{`RANDOM}};
  way0Tag_85 = _RAND_213[20:0];
  _RAND_214 = {1{`RANDOM}};
  way0Tag_86 = _RAND_214[20:0];
  _RAND_215 = {1{`RANDOM}};
  way0Tag_87 = _RAND_215[20:0];
  _RAND_216 = {1{`RANDOM}};
  way0Tag_88 = _RAND_216[20:0];
  _RAND_217 = {1{`RANDOM}};
  way0Tag_89 = _RAND_217[20:0];
  _RAND_218 = {1{`RANDOM}};
  way0Tag_90 = _RAND_218[20:0];
  _RAND_219 = {1{`RANDOM}};
  way0Tag_91 = _RAND_219[20:0];
  _RAND_220 = {1{`RANDOM}};
  way0Tag_92 = _RAND_220[20:0];
  _RAND_221 = {1{`RANDOM}};
  way0Tag_93 = _RAND_221[20:0];
  _RAND_222 = {1{`RANDOM}};
  way0Tag_94 = _RAND_222[20:0];
  _RAND_223 = {1{`RANDOM}};
  way0Tag_95 = _RAND_223[20:0];
  _RAND_224 = {1{`RANDOM}};
  way0Tag_96 = _RAND_224[20:0];
  _RAND_225 = {1{`RANDOM}};
  way0Tag_97 = _RAND_225[20:0];
  _RAND_226 = {1{`RANDOM}};
  way0Tag_98 = _RAND_226[20:0];
  _RAND_227 = {1{`RANDOM}};
  way0Tag_99 = _RAND_227[20:0];
  _RAND_228 = {1{`RANDOM}};
  way0Tag_100 = _RAND_228[20:0];
  _RAND_229 = {1{`RANDOM}};
  way0Tag_101 = _RAND_229[20:0];
  _RAND_230 = {1{`RANDOM}};
  way0Tag_102 = _RAND_230[20:0];
  _RAND_231 = {1{`RANDOM}};
  way0Tag_103 = _RAND_231[20:0];
  _RAND_232 = {1{`RANDOM}};
  way0Tag_104 = _RAND_232[20:0];
  _RAND_233 = {1{`RANDOM}};
  way0Tag_105 = _RAND_233[20:0];
  _RAND_234 = {1{`RANDOM}};
  way0Tag_106 = _RAND_234[20:0];
  _RAND_235 = {1{`RANDOM}};
  way0Tag_107 = _RAND_235[20:0];
  _RAND_236 = {1{`RANDOM}};
  way0Tag_108 = _RAND_236[20:0];
  _RAND_237 = {1{`RANDOM}};
  way0Tag_109 = _RAND_237[20:0];
  _RAND_238 = {1{`RANDOM}};
  way0Tag_110 = _RAND_238[20:0];
  _RAND_239 = {1{`RANDOM}};
  way0Tag_111 = _RAND_239[20:0];
  _RAND_240 = {1{`RANDOM}};
  way0Tag_112 = _RAND_240[20:0];
  _RAND_241 = {1{`RANDOM}};
  way0Tag_113 = _RAND_241[20:0];
  _RAND_242 = {1{`RANDOM}};
  way0Tag_114 = _RAND_242[20:0];
  _RAND_243 = {1{`RANDOM}};
  way0Tag_115 = _RAND_243[20:0];
  _RAND_244 = {1{`RANDOM}};
  way0Tag_116 = _RAND_244[20:0];
  _RAND_245 = {1{`RANDOM}};
  way0Tag_117 = _RAND_245[20:0];
  _RAND_246 = {1{`RANDOM}};
  way0Tag_118 = _RAND_246[20:0];
  _RAND_247 = {1{`RANDOM}};
  way0Tag_119 = _RAND_247[20:0];
  _RAND_248 = {1{`RANDOM}};
  way0Tag_120 = _RAND_248[20:0];
  _RAND_249 = {1{`RANDOM}};
  way0Tag_121 = _RAND_249[20:0];
  _RAND_250 = {1{`RANDOM}};
  way0Tag_122 = _RAND_250[20:0];
  _RAND_251 = {1{`RANDOM}};
  way0Tag_123 = _RAND_251[20:0];
  _RAND_252 = {1{`RANDOM}};
  way0Tag_124 = _RAND_252[20:0];
  _RAND_253 = {1{`RANDOM}};
  way0Tag_125 = _RAND_253[20:0];
  _RAND_254 = {1{`RANDOM}};
  way0Tag_126 = _RAND_254[20:0];
  _RAND_255 = {1{`RANDOM}};
  way0Tag_127 = _RAND_255[20:0];
  _RAND_256 = {1{`RANDOM}};
  way0Age_0 = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  way0Age_1 = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  way0Age_2 = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  way0Age_3 = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  way0Age_4 = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  way0Age_5 = _RAND_261[0:0];
  _RAND_262 = {1{`RANDOM}};
  way0Age_6 = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  way0Age_7 = _RAND_263[0:0];
  _RAND_264 = {1{`RANDOM}};
  way0Age_8 = _RAND_264[0:0];
  _RAND_265 = {1{`RANDOM}};
  way0Age_9 = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  way0Age_10 = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  way0Age_11 = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  way0Age_12 = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  way0Age_13 = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  way0Age_14 = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  way0Age_15 = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  way0Age_16 = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  way0Age_17 = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  way0Age_18 = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  way0Age_19 = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  way0Age_20 = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  way0Age_21 = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  way0Age_22 = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  way0Age_23 = _RAND_279[0:0];
  _RAND_280 = {1{`RANDOM}};
  way0Age_24 = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  way0Age_25 = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  way0Age_26 = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  way0Age_27 = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  way0Age_28 = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  way0Age_29 = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  way0Age_30 = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  way0Age_31 = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  way0Age_32 = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  way0Age_33 = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  way0Age_34 = _RAND_290[0:0];
  _RAND_291 = {1{`RANDOM}};
  way0Age_35 = _RAND_291[0:0];
  _RAND_292 = {1{`RANDOM}};
  way0Age_36 = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  way0Age_37 = _RAND_293[0:0];
  _RAND_294 = {1{`RANDOM}};
  way0Age_38 = _RAND_294[0:0];
  _RAND_295 = {1{`RANDOM}};
  way0Age_39 = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  way0Age_40 = _RAND_296[0:0];
  _RAND_297 = {1{`RANDOM}};
  way0Age_41 = _RAND_297[0:0];
  _RAND_298 = {1{`RANDOM}};
  way0Age_42 = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  way0Age_43 = _RAND_299[0:0];
  _RAND_300 = {1{`RANDOM}};
  way0Age_44 = _RAND_300[0:0];
  _RAND_301 = {1{`RANDOM}};
  way0Age_45 = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  way0Age_46 = _RAND_302[0:0];
  _RAND_303 = {1{`RANDOM}};
  way0Age_47 = _RAND_303[0:0];
  _RAND_304 = {1{`RANDOM}};
  way0Age_48 = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  way0Age_49 = _RAND_305[0:0];
  _RAND_306 = {1{`RANDOM}};
  way0Age_50 = _RAND_306[0:0];
  _RAND_307 = {1{`RANDOM}};
  way0Age_51 = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  way0Age_52 = _RAND_308[0:0];
  _RAND_309 = {1{`RANDOM}};
  way0Age_53 = _RAND_309[0:0];
  _RAND_310 = {1{`RANDOM}};
  way0Age_54 = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  way0Age_55 = _RAND_311[0:0];
  _RAND_312 = {1{`RANDOM}};
  way0Age_56 = _RAND_312[0:0];
  _RAND_313 = {1{`RANDOM}};
  way0Age_57 = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  way0Age_58 = _RAND_314[0:0];
  _RAND_315 = {1{`RANDOM}};
  way0Age_59 = _RAND_315[0:0];
  _RAND_316 = {1{`RANDOM}};
  way0Age_60 = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  way0Age_61 = _RAND_317[0:0];
  _RAND_318 = {1{`RANDOM}};
  way0Age_62 = _RAND_318[0:0];
  _RAND_319 = {1{`RANDOM}};
  way0Age_63 = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  way0Age_64 = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  way0Age_65 = _RAND_321[0:0];
  _RAND_322 = {1{`RANDOM}};
  way0Age_66 = _RAND_322[0:0];
  _RAND_323 = {1{`RANDOM}};
  way0Age_67 = _RAND_323[0:0];
  _RAND_324 = {1{`RANDOM}};
  way0Age_68 = _RAND_324[0:0];
  _RAND_325 = {1{`RANDOM}};
  way0Age_69 = _RAND_325[0:0];
  _RAND_326 = {1{`RANDOM}};
  way0Age_70 = _RAND_326[0:0];
  _RAND_327 = {1{`RANDOM}};
  way0Age_71 = _RAND_327[0:0];
  _RAND_328 = {1{`RANDOM}};
  way0Age_72 = _RAND_328[0:0];
  _RAND_329 = {1{`RANDOM}};
  way0Age_73 = _RAND_329[0:0];
  _RAND_330 = {1{`RANDOM}};
  way0Age_74 = _RAND_330[0:0];
  _RAND_331 = {1{`RANDOM}};
  way0Age_75 = _RAND_331[0:0];
  _RAND_332 = {1{`RANDOM}};
  way0Age_76 = _RAND_332[0:0];
  _RAND_333 = {1{`RANDOM}};
  way0Age_77 = _RAND_333[0:0];
  _RAND_334 = {1{`RANDOM}};
  way0Age_78 = _RAND_334[0:0];
  _RAND_335 = {1{`RANDOM}};
  way0Age_79 = _RAND_335[0:0];
  _RAND_336 = {1{`RANDOM}};
  way0Age_80 = _RAND_336[0:0];
  _RAND_337 = {1{`RANDOM}};
  way0Age_81 = _RAND_337[0:0];
  _RAND_338 = {1{`RANDOM}};
  way0Age_82 = _RAND_338[0:0];
  _RAND_339 = {1{`RANDOM}};
  way0Age_83 = _RAND_339[0:0];
  _RAND_340 = {1{`RANDOM}};
  way0Age_84 = _RAND_340[0:0];
  _RAND_341 = {1{`RANDOM}};
  way0Age_85 = _RAND_341[0:0];
  _RAND_342 = {1{`RANDOM}};
  way0Age_86 = _RAND_342[0:0];
  _RAND_343 = {1{`RANDOM}};
  way0Age_87 = _RAND_343[0:0];
  _RAND_344 = {1{`RANDOM}};
  way0Age_88 = _RAND_344[0:0];
  _RAND_345 = {1{`RANDOM}};
  way0Age_89 = _RAND_345[0:0];
  _RAND_346 = {1{`RANDOM}};
  way0Age_90 = _RAND_346[0:0];
  _RAND_347 = {1{`RANDOM}};
  way0Age_91 = _RAND_347[0:0];
  _RAND_348 = {1{`RANDOM}};
  way0Age_92 = _RAND_348[0:0];
  _RAND_349 = {1{`RANDOM}};
  way0Age_93 = _RAND_349[0:0];
  _RAND_350 = {1{`RANDOM}};
  way0Age_94 = _RAND_350[0:0];
  _RAND_351 = {1{`RANDOM}};
  way0Age_95 = _RAND_351[0:0];
  _RAND_352 = {1{`RANDOM}};
  way0Age_96 = _RAND_352[0:0];
  _RAND_353 = {1{`RANDOM}};
  way0Age_97 = _RAND_353[0:0];
  _RAND_354 = {1{`RANDOM}};
  way0Age_98 = _RAND_354[0:0];
  _RAND_355 = {1{`RANDOM}};
  way0Age_99 = _RAND_355[0:0];
  _RAND_356 = {1{`RANDOM}};
  way0Age_100 = _RAND_356[0:0];
  _RAND_357 = {1{`RANDOM}};
  way0Age_101 = _RAND_357[0:0];
  _RAND_358 = {1{`RANDOM}};
  way0Age_102 = _RAND_358[0:0];
  _RAND_359 = {1{`RANDOM}};
  way0Age_103 = _RAND_359[0:0];
  _RAND_360 = {1{`RANDOM}};
  way0Age_104 = _RAND_360[0:0];
  _RAND_361 = {1{`RANDOM}};
  way0Age_105 = _RAND_361[0:0];
  _RAND_362 = {1{`RANDOM}};
  way0Age_106 = _RAND_362[0:0];
  _RAND_363 = {1{`RANDOM}};
  way0Age_107 = _RAND_363[0:0];
  _RAND_364 = {1{`RANDOM}};
  way0Age_108 = _RAND_364[0:0];
  _RAND_365 = {1{`RANDOM}};
  way0Age_109 = _RAND_365[0:0];
  _RAND_366 = {1{`RANDOM}};
  way0Age_110 = _RAND_366[0:0];
  _RAND_367 = {1{`RANDOM}};
  way0Age_111 = _RAND_367[0:0];
  _RAND_368 = {1{`RANDOM}};
  way0Age_112 = _RAND_368[0:0];
  _RAND_369 = {1{`RANDOM}};
  way0Age_113 = _RAND_369[0:0];
  _RAND_370 = {1{`RANDOM}};
  way0Age_114 = _RAND_370[0:0];
  _RAND_371 = {1{`RANDOM}};
  way0Age_115 = _RAND_371[0:0];
  _RAND_372 = {1{`RANDOM}};
  way0Age_116 = _RAND_372[0:0];
  _RAND_373 = {1{`RANDOM}};
  way0Age_117 = _RAND_373[0:0];
  _RAND_374 = {1{`RANDOM}};
  way0Age_118 = _RAND_374[0:0];
  _RAND_375 = {1{`RANDOM}};
  way0Age_119 = _RAND_375[0:0];
  _RAND_376 = {1{`RANDOM}};
  way0Age_120 = _RAND_376[0:0];
  _RAND_377 = {1{`RANDOM}};
  way0Age_121 = _RAND_377[0:0];
  _RAND_378 = {1{`RANDOM}};
  way0Age_122 = _RAND_378[0:0];
  _RAND_379 = {1{`RANDOM}};
  way0Age_123 = _RAND_379[0:0];
  _RAND_380 = {1{`RANDOM}};
  way0Age_124 = _RAND_380[0:0];
  _RAND_381 = {1{`RANDOM}};
  way0Age_125 = _RAND_381[0:0];
  _RAND_382 = {1{`RANDOM}};
  way0Age_126 = _RAND_382[0:0];
  _RAND_383 = {1{`RANDOM}};
  way0Age_127 = _RAND_383[0:0];
  _RAND_384 = {1{`RANDOM}};
  way0Dirty_0 = _RAND_384[0:0];
  _RAND_385 = {1{`RANDOM}};
  way0Dirty_1 = _RAND_385[0:0];
  _RAND_386 = {1{`RANDOM}};
  way0Dirty_2 = _RAND_386[0:0];
  _RAND_387 = {1{`RANDOM}};
  way0Dirty_3 = _RAND_387[0:0];
  _RAND_388 = {1{`RANDOM}};
  way0Dirty_4 = _RAND_388[0:0];
  _RAND_389 = {1{`RANDOM}};
  way0Dirty_5 = _RAND_389[0:0];
  _RAND_390 = {1{`RANDOM}};
  way0Dirty_6 = _RAND_390[0:0];
  _RAND_391 = {1{`RANDOM}};
  way0Dirty_7 = _RAND_391[0:0];
  _RAND_392 = {1{`RANDOM}};
  way0Dirty_8 = _RAND_392[0:0];
  _RAND_393 = {1{`RANDOM}};
  way0Dirty_9 = _RAND_393[0:0];
  _RAND_394 = {1{`RANDOM}};
  way0Dirty_10 = _RAND_394[0:0];
  _RAND_395 = {1{`RANDOM}};
  way0Dirty_11 = _RAND_395[0:0];
  _RAND_396 = {1{`RANDOM}};
  way0Dirty_12 = _RAND_396[0:0];
  _RAND_397 = {1{`RANDOM}};
  way0Dirty_13 = _RAND_397[0:0];
  _RAND_398 = {1{`RANDOM}};
  way0Dirty_14 = _RAND_398[0:0];
  _RAND_399 = {1{`RANDOM}};
  way0Dirty_15 = _RAND_399[0:0];
  _RAND_400 = {1{`RANDOM}};
  way0Dirty_16 = _RAND_400[0:0];
  _RAND_401 = {1{`RANDOM}};
  way0Dirty_17 = _RAND_401[0:0];
  _RAND_402 = {1{`RANDOM}};
  way0Dirty_18 = _RAND_402[0:0];
  _RAND_403 = {1{`RANDOM}};
  way0Dirty_19 = _RAND_403[0:0];
  _RAND_404 = {1{`RANDOM}};
  way0Dirty_20 = _RAND_404[0:0];
  _RAND_405 = {1{`RANDOM}};
  way0Dirty_21 = _RAND_405[0:0];
  _RAND_406 = {1{`RANDOM}};
  way0Dirty_22 = _RAND_406[0:0];
  _RAND_407 = {1{`RANDOM}};
  way0Dirty_23 = _RAND_407[0:0];
  _RAND_408 = {1{`RANDOM}};
  way0Dirty_24 = _RAND_408[0:0];
  _RAND_409 = {1{`RANDOM}};
  way0Dirty_25 = _RAND_409[0:0];
  _RAND_410 = {1{`RANDOM}};
  way0Dirty_26 = _RAND_410[0:0];
  _RAND_411 = {1{`RANDOM}};
  way0Dirty_27 = _RAND_411[0:0];
  _RAND_412 = {1{`RANDOM}};
  way0Dirty_28 = _RAND_412[0:0];
  _RAND_413 = {1{`RANDOM}};
  way0Dirty_29 = _RAND_413[0:0];
  _RAND_414 = {1{`RANDOM}};
  way0Dirty_30 = _RAND_414[0:0];
  _RAND_415 = {1{`RANDOM}};
  way0Dirty_31 = _RAND_415[0:0];
  _RAND_416 = {1{`RANDOM}};
  way0Dirty_32 = _RAND_416[0:0];
  _RAND_417 = {1{`RANDOM}};
  way0Dirty_33 = _RAND_417[0:0];
  _RAND_418 = {1{`RANDOM}};
  way0Dirty_34 = _RAND_418[0:0];
  _RAND_419 = {1{`RANDOM}};
  way0Dirty_35 = _RAND_419[0:0];
  _RAND_420 = {1{`RANDOM}};
  way0Dirty_36 = _RAND_420[0:0];
  _RAND_421 = {1{`RANDOM}};
  way0Dirty_37 = _RAND_421[0:0];
  _RAND_422 = {1{`RANDOM}};
  way0Dirty_38 = _RAND_422[0:0];
  _RAND_423 = {1{`RANDOM}};
  way0Dirty_39 = _RAND_423[0:0];
  _RAND_424 = {1{`RANDOM}};
  way0Dirty_40 = _RAND_424[0:0];
  _RAND_425 = {1{`RANDOM}};
  way0Dirty_41 = _RAND_425[0:0];
  _RAND_426 = {1{`RANDOM}};
  way0Dirty_42 = _RAND_426[0:0];
  _RAND_427 = {1{`RANDOM}};
  way0Dirty_43 = _RAND_427[0:0];
  _RAND_428 = {1{`RANDOM}};
  way0Dirty_44 = _RAND_428[0:0];
  _RAND_429 = {1{`RANDOM}};
  way0Dirty_45 = _RAND_429[0:0];
  _RAND_430 = {1{`RANDOM}};
  way0Dirty_46 = _RAND_430[0:0];
  _RAND_431 = {1{`RANDOM}};
  way0Dirty_47 = _RAND_431[0:0];
  _RAND_432 = {1{`RANDOM}};
  way0Dirty_48 = _RAND_432[0:0];
  _RAND_433 = {1{`RANDOM}};
  way0Dirty_49 = _RAND_433[0:0];
  _RAND_434 = {1{`RANDOM}};
  way0Dirty_50 = _RAND_434[0:0];
  _RAND_435 = {1{`RANDOM}};
  way0Dirty_51 = _RAND_435[0:0];
  _RAND_436 = {1{`RANDOM}};
  way0Dirty_52 = _RAND_436[0:0];
  _RAND_437 = {1{`RANDOM}};
  way0Dirty_53 = _RAND_437[0:0];
  _RAND_438 = {1{`RANDOM}};
  way0Dirty_54 = _RAND_438[0:0];
  _RAND_439 = {1{`RANDOM}};
  way0Dirty_55 = _RAND_439[0:0];
  _RAND_440 = {1{`RANDOM}};
  way0Dirty_56 = _RAND_440[0:0];
  _RAND_441 = {1{`RANDOM}};
  way0Dirty_57 = _RAND_441[0:0];
  _RAND_442 = {1{`RANDOM}};
  way0Dirty_58 = _RAND_442[0:0];
  _RAND_443 = {1{`RANDOM}};
  way0Dirty_59 = _RAND_443[0:0];
  _RAND_444 = {1{`RANDOM}};
  way0Dirty_60 = _RAND_444[0:0];
  _RAND_445 = {1{`RANDOM}};
  way0Dirty_61 = _RAND_445[0:0];
  _RAND_446 = {1{`RANDOM}};
  way0Dirty_62 = _RAND_446[0:0];
  _RAND_447 = {1{`RANDOM}};
  way0Dirty_63 = _RAND_447[0:0];
  _RAND_448 = {1{`RANDOM}};
  way0Dirty_64 = _RAND_448[0:0];
  _RAND_449 = {1{`RANDOM}};
  way0Dirty_65 = _RAND_449[0:0];
  _RAND_450 = {1{`RANDOM}};
  way0Dirty_66 = _RAND_450[0:0];
  _RAND_451 = {1{`RANDOM}};
  way0Dirty_67 = _RAND_451[0:0];
  _RAND_452 = {1{`RANDOM}};
  way0Dirty_68 = _RAND_452[0:0];
  _RAND_453 = {1{`RANDOM}};
  way0Dirty_69 = _RAND_453[0:0];
  _RAND_454 = {1{`RANDOM}};
  way0Dirty_70 = _RAND_454[0:0];
  _RAND_455 = {1{`RANDOM}};
  way0Dirty_71 = _RAND_455[0:0];
  _RAND_456 = {1{`RANDOM}};
  way0Dirty_72 = _RAND_456[0:0];
  _RAND_457 = {1{`RANDOM}};
  way0Dirty_73 = _RAND_457[0:0];
  _RAND_458 = {1{`RANDOM}};
  way0Dirty_74 = _RAND_458[0:0];
  _RAND_459 = {1{`RANDOM}};
  way0Dirty_75 = _RAND_459[0:0];
  _RAND_460 = {1{`RANDOM}};
  way0Dirty_76 = _RAND_460[0:0];
  _RAND_461 = {1{`RANDOM}};
  way0Dirty_77 = _RAND_461[0:0];
  _RAND_462 = {1{`RANDOM}};
  way0Dirty_78 = _RAND_462[0:0];
  _RAND_463 = {1{`RANDOM}};
  way0Dirty_79 = _RAND_463[0:0];
  _RAND_464 = {1{`RANDOM}};
  way0Dirty_80 = _RAND_464[0:0];
  _RAND_465 = {1{`RANDOM}};
  way0Dirty_81 = _RAND_465[0:0];
  _RAND_466 = {1{`RANDOM}};
  way0Dirty_82 = _RAND_466[0:0];
  _RAND_467 = {1{`RANDOM}};
  way0Dirty_83 = _RAND_467[0:0];
  _RAND_468 = {1{`RANDOM}};
  way0Dirty_84 = _RAND_468[0:0];
  _RAND_469 = {1{`RANDOM}};
  way0Dirty_85 = _RAND_469[0:0];
  _RAND_470 = {1{`RANDOM}};
  way0Dirty_86 = _RAND_470[0:0];
  _RAND_471 = {1{`RANDOM}};
  way0Dirty_87 = _RAND_471[0:0];
  _RAND_472 = {1{`RANDOM}};
  way0Dirty_88 = _RAND_472[0:0];
  _RAND_473 = {1{`RANDOM}};
  way0Dirty_89 = _RAND_473[0:0];
  _RAND_474 = {1{`RANDOM}};
  way0Dirty_90 = _RAND_474[0:0];
  _RAND_475 = {1{`RANDOM}};
  way0Dirty_91 = _RAND_475[0:0];
  _RAND_476 = {1{`RANDOM}};
  way0Dirty_92 = _RAND_476[0:0];
  _RAND_477 = {1{`RANDOM}};
  way0Dirty_93 = _RAND_477[0:0];
  _RAND_478 = {1{`RANDOM}};
  way0Dirty_94 = _RAND_478[0:0];
  _RAND_479 = {1{`RANDOM}};
  way0Dirty_95 = _RAND_479[0:0];
  _RAND_480 = {1{`RANDOM}};
  way0Dirty_96 = _RAND_480[0:0];
  _RAND_481 = {1{`RANDOM}};
  way0Dirty_97 = _RAND_481[0:0];
  _RAND_482 = {1{`RANDOM}};
  way0Dirty_98 = _RAND_482[0:0];
  _RAND_483 = {1{`RANDOM}};
  way0Dirty_99 = _RAND_483[0:0];
  _RAND_484 = {1{`RANDOM}};
  way0Dirty_100 = _RAND_484[0:0];
  _RAND_485 = {1{`RANDOM}};
  way0Dirty_101 = _RAND_485[0:0];
  _RAND_486 = {1{`RANDOM}};
  way0Dirty_102 = _RAND_486[0:0];
  _RAND_487 = {1{`RANDOM}};
  way0Dirty_103 = _RAND_487[0:0];
  _RAND_488 = {1{`RANDOM}};
  way0Dirty_104 = _RAND_488[0:0];
  _RAND_489 = {1{`RANDOM}};
  way0Dirty_105 = _RAND_489[0:0];
  _RAND_490 = {1{`RANDOM}};
  way0Dirty_106 = _RAND_490[0:0];
  _RAND_491 = {1{`RANDOM}};
  way0Dirty_107 = _RAND_491[0:0];
  _RAND_492 = {1{`RANDOM}};
  way0Dirty_108 = _RAND_492[0:0];
  _RAND_493 = {1{`RANDOM}};
  way0Dirty_109 = _RAND_493[0:0];
  _RAND_494 = {1{`RANDOM}};
  way0Dirty_110 = _RAND_494[0:0];
  _RAND_495 = {1{`RANDOM}};
  way0Dirty_111 = _RAND_495[0:0];
  _RAND_496 = {1{`RANDOM}};
  way0Dirty_112 = _RAND_496[0:0];
  _RAND_497 = {1{`RANDOM}};
  way0Dirty_113 = _RAND_497[0:0];
  _RAND_498 = {1{`RANDOM}};
  way0Dirty_114 = _RAND_498[0:0];
  _RAND_499 = {1{`RANDOM}};
  way0Dirty_115 = _RAND_499[0:0];
  _RAND_500 = {1{`RANDOM}};
  way0Dirty_116 = _RAND_500[0:0];
  _RAND_501 = {1{`RANDOM}};
  way0Dirty_117 = _RAND_501[0:0];
  _RAND_502 = {1{`RANDOM}};
  way0Dirty_118 = _RAND_502[0:0];
  _RAND_503 = {1{`RANDOM}};
  way0Dirty_119 = _RAND_503[0:0];
  _RAND_504 = {1{`RANDOM}};
  way0Dirty_120 = _RAND_504[0:0];
  _RAND_505 = {1{`RANDOM}};
  way0Dirty_121 = _RAND_505[0:0];
  _RAND_506 = {1{`RANDOM}};
  way0Dirty_122 = _RAND_506[0:0];
  _RAND_507 = {1{`RANDOM}};
  way0Dirty_123 = _RAND_507[0:0];
  _RAND_508 = {1{`RANDOM}};
  way0Dirty_124 = _RAND_508[0:0];
  _RAND_509 = {1{`RANDOM}};
  way0Dirty_125 = _RAND_509[0:0];
  _RAND_510 = {1{`RANDOM}};
  way0Dirty_126 = _RAND_510[0:0];
  _RAND_511 = {1{`RANDOM}};
  way0Dirty_127 = _RAND_511[0:0];
  _RAND_512 = {1{`RANDOM}};
  way1V_0 = _RAND_512[0:0];
  _RAND_513 = {1{`RANDOM}};
  way1V_1 = _RAND_513[0:0];
  _RAND_514 = {1{`RANDOM}};
  way1V_2 = _RAND_514[0:0];
  _RAND_515 = {1{`RANDOM}};
  way1V_3 = _RAND_515[0:0];
  _RAND_516 = {1{`RANDOM}};
  way1V_4 = _RAND_516[0:0];
  _RAND_517 = {1{`RANDOM}};
  way1V_5 = _RAND_517[0:0];
  _RAND_518 = {1{`RANDOM}};
  way1V_6 = _RAND_518[0:0];
  _RAND_519 = {1{`RANDOM}};
  way1V_7 = _RAND_519[0:0];
  _RAND_520 = {1{`RANDOM}};
  way1V_8 = _RAND_520[0:0];
  _RAND_521 = {1{`RANDOM}};
  way1V_9 = _RAND_521[0:0];
  _RAND_522 = {1{`RANDOM}};
  way1V_10 = _RAND_522[0:0];
  _RAND_523 = {1{`RANDOM}};
  way1V_11 = _RAND_523[0:0];
  _RAND_524 = {1{`RANDOM}};
  way1V_12 = _RAND_524[0:0];
  _RAND_525 = {1{`RANDOM}};
  way1V_13 = _RAND_525[0:0];
  _RAND_526 = {1{`RANDOM}};
  way1V_14 = _RAND_526[0:0];
  _RAND_527 = {1{`RANDOM}};
  way1V_15 = _RAND_527[0:0];
  _RAND_528 = {1{`RANDOM}};
  way1V_16 = _RAND_528[0:0];
  _RAND_529 = {1{`RANDOM}};
  way1V_17 = _RAND_529[0:0];
  _RAND_530 = {1{`RANDOM}};
  way1V_18 = _RAND_530[0:0];
  _RAND_531 = {1{`RANDOM}};
  way1V_19 = _RAND_531[0:0];
  _RAND_532 = {1{`RANDOM}};
  way1V_20 = _RAND_532[0:0];
  _RAND_533 = {1{`RANDOM}};
  way1V_21 = _RAND_533[0:0];
  _RAND_534 = {1{`RANDOM}};
  way1V_22 = _RAND_534[0:0];
  _RAND_535 = {1{`RANDOM}};
  way1V_23 = _RAND_535[0:0];
  _RAND_536 = {1{`RANDOM}};
  way1V_24 = _RAND_536[0:0];
  _RAND_537 = {1{`RANDOM}};
  way1V_25 = _RAND_537[0:0];
  _RAND_538 = {1{`RANDOM}};
  way1V_26 = _RAND_538[0:0];
  _RAND_539 = {1{`RANDOM}};
  way1V_27 = _RAND_539[0:0];
  _RAND_540 = {1{`RANDOM}};
  way1V_28 = _RAND_540[0:0];
  _RAND_541 = {1{`RANDOM}};
  way1V_29 = _RAND_541[0:0];
  _RAND_542 = {1{`RANDOM}};
  way1V_30 = _RAND_542[0:0];
  _RAND_543 = {1{`RANDOM}};
  way1V_31 = _RAND_543[0:0];
  _RAND_544 = {1{`RANDOM}};
  way1V_32 = _RAND_544[0:0];
  _RAND_545 = {1{`RANDOM}};
  way1V_33 = _RAND_545[0:0];
  _RAND_546 = {1{`RANDOM}};
  way1V_34 = _RAND_546[0:0];
  _RAND_547 = {1{`RANDOM}};
  way1V_35 = _RAND_547[0:0];
  _RAND_548 = {1{`RANDOM}};
  way1V_36 = _RAND_548[0:0];
  _RAND_549 = {1{`RANDOM}};
  way1V_37 = _RAND_549[0:0];
  _RAND_550 = {1{`RANDOM}};
  way1V_38 = _RAND_550[0:0];
  _RAND_551 = {1{`RANDOM}};
  way1V_39 = _RAND_551[0:0];
  _RAND_552 = {1{`RANDOM}};
  way1V_40 = _RAND_552[0:0];
  _RAND_553 = {1{`RANDOM}};
  way1V_41 = _RAND_553[0:0];
  _RAND_554 = {1{`RANDOM}};
  way1V_42 = _RAND_554[0:0];
  _RAND_555 = {1{`RANDOM}};
  way1V_43 = _RAND_555[0:0];
  _RAND_556 = {1{`RANDOM}};
  way1V_44 = _RAND_556[0:0];
  _RAND_557 = {1{`RANDOM}};
  way1V_45 = _RAND_557[0:0];
  _RAND_558 = {1{`RANDOM}};
  way1V_46 = _RAND_558[0:0];
  _RAND_559 = {1{`RANDOM}};
  way1V_47 = _RAND_559[0:0];
  _RAND_560 = {1{`RANDOM}};
  way1V_48 = _RAND_560[0:0];
  _RAND_561 = {1{`RANDOM}};
  way1V_49 = _RAND_561[0:0];
  _RAND_562 = {1{`RANDOM}};
  way1V_50 = _RAND_562[0:0];
  _RAND_563 = {1{`RANDOM}};
  way1V_51 = _RAND_563[0:0];
  _RAND_564 = {1{`RANDOM}};
  way1V_52 = _RAND_564[0:0];
  _RAND_565 = {1{`RANDOM}};
  way1V_53 = _RAND_565[0:0];
  _RAND_566 = {1{`RANDOM}};
  way1V_54 = _RAND_566[0:0];
  _RAND_567 = {1{`RANDOM}};
  way1V_55 = _RAND_567[0:0];
  _RAND_568 = {1{`RANDOM}};
  way1V_56 = _RAND_568[0:0];
  _RAND_569 = {1{`RANDOM}};
  way1V_57 = _RAND_569[0:0];
  _RAND_570 = {1{`RANDOM}};
  way1V_58 = _RAND_570[0:0];
  _RAND_571 = {1{`RANDOM}};
  way1V_59 = _RAND_571[0:0];
  _RAND_572 = {1{`RANDOM}};
  way1V_60 = _RAND_572[0:0];
  _RAND_573 = {1{`RANDOM}};
  way1V_61 = _RAND_573[0:0];
  _RAND_574 = {1{`RANDOM}};
  way1V_62 = _RAND_574[0:0];
  _RAND_575 = {1{`RANDOM}};
  way1V_63 = _RAND_575[0:0];
  _RAND_576 = {1{`RANDOM}};
  way1V_64 = _RAND_576[0:0];
  _RAND_577 = {1{`RANDOM}};
  way1V_65 = _RAND_577[0:0];
  _RAND_578 = {1{`RANDOM}};
  way1V_66 = _RAND_578[0:0];
  _RAND_579 = {1{`RANDOM}};
  way1V_67 = _RAND_579[0:0];
  _RAND_580 = {1{`RANDOM}};
  way1V_68 = _RAND_580[0:0];
  _RAND_581 = {1{`RANDOM}};
  way1V_69 = _RAND_581[0:0];
  _RAND_582 = {1{`RANDOM}};
  way1V_70 = _RAND_582[0:0];
  _RAND_583 = {1{`RANDOM}};
  way1V_71 = _RAND_583[0:0];
  _RAND_584 = {1{`RANDOM}};
  way1V_72 = _RAND_584[0:0];
  _RAND_585 = {1{`RANDOM}};
  way1V_73 = _RAND_585[0:0];
  _RAND_586 = {1{`RANDOM}};
  way1V_74 = _RAND_586[0:0];
  _RAND_587 = {1{`RANDOM}};
  way1V_75 = _RAND_587[0:0];
  _RAND_588 = {1{`RANDOM}};
  way1V_76 = _RAND_588[0:0];
  _RAND_589 = {1{`RANDOM}};
  way1V_77 = _RAND_589[0:0];
  _RAND_590 = {1{`RANDOM}};
  way1V_78 = _RAND_590[0:0];
  _RAND_591 = {1{`RANDOM}};
  way1V_79 = _RAND_591[0:0];
  _RAND_592 = {1{`RANDOM}};
  way1V_80 = _RAND_592[0:0];
  _RAND_593 = {1{`RANDOM}};
  way1V_81 = _RAND_593[0:0];
  _RAND_594 = {1{`RANDOM}};
  way1V_82 = _RAND_594[0:0];
  _RAND_595 = {1{`RANDOM}};
  way1V_83 = _RAND_595[0:0];
  _RAND_596 = {1{`RANDOM}};
  way1V_84 = _RAND_596[0:0];
  _RAND_597 = {1{`RANDOM}};
  way1V_85 = _RAND_597[0:0];
  _RAND_598 = {1{`RANDOM}};
  way1V_86 = _RAND_598[0:0];
  _RAND_599 = {1{`RANDOM}};
  way1V_87 = _RAND_599[0:0];
  _RAND_600 = {1{`RANDOM}};
  way1V_88 = _RAND_600[0:0];
  _RAND_601 = {1{`RANDOM}};
  way1V_89 = _RAND_601[0:0];
  _RAND_602 = {1{`RANDOM}};
  way1V_90 = _RAND_602[0:0];
  _RAND_603 = {1{`RANDOM}};
  way1V_91 = _RAND_603[0:0];
  _RAND_604 = {1{`RANDOM}};
  way1V_92 = _RAND_604[0:0];
  _RAND_605 = {1{`RANDOM}};
  way1V_93 = _RAND_605[0:0];
  _RAND_606 = {1{`RANDOM}};
  way1V_94 = _RAND_606[0:0];
  _RAND_607 = {1{`RANDOM}};
  way1V_95 = _RAND_607[0:0];
  _RAND_608 = {1{`RANDOM}};
  way1V_96 = _RAND_608[0:0];
  _RAND_609 = {1{`RANDOM}};
  way1V_97 = _RAND_609[0:0];
  _RAND_610 = {1{`RANDOM}};
  way1V_98 = _RAND_610[0:0];
  _RAND_611 = {1{`RANDOM}};
  way1V_99 = _RAND_611[0:0];
  _RAND_612 = {1{`RANDOM}};
  way1V_100 = _RAND_612[0:0];
  _RAND_613 = {1{`RANDOM}};
  way1V_101 = _RAND_613[0:0];
  _RAND_614 = {1{`RANDOM}};
  way1V_102 = _RAND_614[0:0];
  _RAND_615 = {1{`RANDOM}};
  way1V_103 = _RAND_615[0:0];
  _RAND_616 = {1{`RANDOM}};
  way1V_104 = _RAND_616[0:0];
  _RAND_617 = {1{`RANDOM}};
  way1V_105 = _RAND_617[0:0];
  _RAND_618 = {1{`RANDOM}};
  way1V_106 = _RAND_618[0:0];
  _RAND_619 = {1{`RANDOM}};
  way1V_107 = _RAND_619[0:0];
  _RAND_620 = {1{`RANDOM}};
  way1V_108 = _RAND_620[0:0];
  _RAND_621 = {1{`RANDOM}};
  way1V_109 = _RAND_621[0:0];
  _RAND_622 = {1{`RANDOM}};
  way1V_110 = _RAND_622[0:0];
  _RAND_623 = {1{`RANDOM}};
  way1V_111 = _RAND_623[0:0];
  _RAND_624 = {1{`RANDOM}};
  way1V_112 = _RAND_624[0:0];
  _RAND_625 = {1{`RANDOM}};
  way1V_113 = _RAND_625[0:0];
  _RAND_626 = {1{`RANDOM}};
  way1V_114 = _RAND_626[0:0];
  _RAND_627 = {1{`RANDOM}};
  way1V_115 = _RAND_627[0:0];
  _RAND_628 = {1{`RANDOM}};
  way1V_116 = _RAND_628[0:0];
  _RAND_629 = {1{`RANDOM}};
  way1V_117 = _RAND_629[0:0];
  _RAND_630 = {1{`RANDOM}};
  way1V_118 = _RAND_630[0:0];
  _RAND_631 = {1{`RANDOM}};
  way1V_119 = _RAND_631[0:0];
  _RAND_632 = {1{`RANDOM}};
  way1V_120 = _RAND_632[0:0];
  _RAND_633 = {1{`RANDOM}};
  way1V_121 = _RAND_633[0:0];
  _RAND_634 = {1{`RANDOM}};
  way1V_122 = _RAND_634[0:0];
  _RAND_635 = {1{`RANDOM}};
  way1V_123 = _RAND_635[0:0];
  _RAND_636 = {1{`RANDOM}};
  way1V_124 = _RAND_636[0:0];
  _RAND_637 = {1{`RANDOM}};
  way1V_125 = _RAND_637[0:0];
  _RAND_638 = {1{`RANDOM}};
  way1V_126 = _RAND_638[0:0];
  _RAND_639 = {1{`RANDOM}};
  way1V_127 = _RAND_639[0:0];
  _RAND_640 = {1{`RANDOM}};
  way1Tag_0 = _RAND_640[20:0];
  _RAND_641 = {1{`RANDOM}};
  way1Tag_1 = _RAND_641[20:0];
  _RAND_642 = {1{`RANDOM}};
  way1Tag_2 = _RAND_642[20:0];
  _RAND_643 = {1{`RANDOM}};
  way1Tag_3 = _RAND_643[20:0];
  _RAND_644 = {1{`RANDOM}};
  way1Tag_4 = _RAND_644[20:0];
  _RAND_645 = {1{`RANDOM}};
  way1Tag_5 = _RAND_645[20:0];
  _RAND_646 = {1{`RANDOM}};
  way1Tag_6 = _RAND_646[20:0];
  _RAND_647 = {1{`RANDOM}};
  way1Tag_7 = _RAND_647[20:0];
  _RAND_648 = {1{`RANDOM}};
  way1Tag_8 = _RAND_648[20:0];
  _RAND_649 = {1{`RANDOM}};
  way1Tag_9 = _RAND_649[20:0];
  _RAND_650 = {1{`RANDOM}};
  way1Tag_10 = _RAND_650[20:0];
  _RAND_651 = {1{`RANDOM}};
  way1Tag_11 = _RAND_651[20:0];
  _RAND_652 = {1{`RANDOM}};
  way1Tag_12 = _RAND_652[20:0];
  _RAND_653 = {1{`RANDOM}};
  way1Tag_13 = _RAND_653[20:0];
  _RAND_654 = {1{`RANDOM}};
  way1Tag_14 = _RAND_654[20:0];
  _RAND_655 = {1{`RANDOM}};
  way1Tag_15 = _RAND_655[20:0];
  _RAND_656 = {1{`RANDOM}};
  way1Tag_16 = _RAND_656[20:0];
  _RAND_657 = {1{`RANDOM}};
  way1Tag_17 = _RAND_657[20:0];
  _RAND_658 = {1{`RANDOM}};
  way1Tag_18 = _RAND_658[20:0];
  _RAND_659 = {1{`RANDOM}};
  way1Tag_19 = _RAND_659[20:0];
  _RAND_660 = {1{`RANDOM}};
  way1Tag_20 = _RAND_660[20:0];
  _RAND_661 = {1{`RANDOM}};
  way1Tag_21 = _RAND_661[20:0];
  _RAND_662 = {1{`RANDOM}};
  way1Tag_22 = _RAND_662[20:0];
  _RAND_663 = {1{`RANDOM}};
  way1Tag_23 = _RAND_663[20:0];
  _RAND_664 = {1{`RANDOM}};
  way1Tag_24 = _RAND_664[20:0];
  _RAND_665 = {1{`RANDOM}};
  way1Tag_25 = _RAND_665[20:0];
  _RAND_666 = {1{`RANDOM}};
  way1Tag_26 = _RAND_666[20:0];
  _RAND_667 = {1{`RANDOM}};
  way1Tag_27 = _RAND_667[20:0];
  _RAND_668 = {1{`RANDOM}};
  way1Tag_28 = _RAND_668[20:0];
  _RAND_669 = {1{`RANDOM}};
  way1Tag_29 = _RAND_669[20:0];
  _RAND_670 = {1{`RANDOM}};
  way1Tag_30 = _RAND_670[20:0];
  _RAND_671 = {1{`RANDOM}};
  way1Tag_31 = _RAND_671[20:0];
  _RAND_672 = {1{`RANDOM}};
  way1Tag_32 = _RAND_672[20:0];
  _RAND_673 = {1{`RANDOM}};
  way1Tag_33 = _RAND_673[20:0];
  _RAND_674 = {1{`RANDOM}};
  way1Tag_34 = _RAND_674[20:0];
  _RAND_675 = {1{`RANDOM}};
  way1Tag_35 = _RAND_675[20:0];
  _RAND_676 = {1{`RANDOM}};
  way1Tag_36 = _RAND_676[20:0];
  _RAND_677 = {1{`RANDOM}};
  way1Tag_37 = _RAND_677[20:0];
  _RAND_678 = {1{`RANDOM}};
  way1Tag_38 = _RAND_678[20:0];
  _RAND_679 = {1{`RANDOM}};
  way1Tag_39 = _RAND_679[20:0];
  _RAND_680 = {1{`RANDOM}};
  way1Tag_40 = _RAND_680[20:0];
  _RAND_681 = {1{`RANDOM}};
  way1Tag_41 = _RAND_681[20:0];
  _RAND_682 = {1{`RANDOM}};
  way1Tag_42 = _RAND_682[20:0];
  _RAND_683 = {1{`RANDOM}};
  way1Tag_43 = _RAND_683[20:0];
  _RAND_684 = {1{`RANDOM}};
  way1Tag_44 = _RAND_684[20:0];
  _RAND_685 = {1{`RANDOM}};
  way1Tag_45 = _RAND_685[20:0];
  _RAND_686 = {1{`RANDOM}};
  way1Tag_46 = _RAND_686[20:0];
  _RAND_687 = {1{`RANDOM}};
  way1Tag_47 = _RAND_687[20:0];
  _RAND_688 = {1{`RANDOM}};
  way1Tag_48 = _RAND_688[20:0];
  _RAND_689 = {1{`RANDOM}};
  way1Tag_49 = _RAND_689[20:0];
  _RAND_690 = {1{`RANDOM}};
  way1Tag_50 = _RAND_690[20:0];
  _RAND_691 = {1{`RANDOM}};
  way1Tag_51 = _RAND_691[20:0];
  _RAND_692 = {1{`RANDOM}};
  way1Tag_52 = _RAND_692[20:0];
  _RAND_693 = {1{`RANDOM}};
  way1Tag_53 = _RAND_693[20:0];
  _RAND_694 = {1{`RANDOM}};
  way1Tag_54 = _RAND_694[20:0];
  _RAND_695 = {1{`RANDOM}};
  way1Tag_55 = _RAND_695[20:0];
  _RAND_696 = {1{`RANDOM}};
  way1Tag_56 = _RAND_696[20:0];
  _RAND_697 = {1{`RANDOM}};
  way1Tag_57 = _RAND_697[20:0];
  _RAND_698 = {1{`RANDOM}};
  way1Tag_58 = _RAND_698[20:0];
  _RAND_699 = {1{`RANDOM}};
  way1Tag_59 = _RAND_699[20:0];
  _RAND_700 = {1{`RANDOM}};
  way1Tag_60 = _RAND_700[20:0];
  _RAND_701 = {1{`RANDOM}};
  way1Tag_61 = _RAND_701[20:0];
  _RAND_702 = {1{`RANDOM}};
  way1Tag_62 = _RAND_702[20:0];
  _RAND_703 = {1{`RANDOM}};
  way1Tag_63 = _RAND_703[20:0];
  _RAND_704 = {1{`RANDOM}};
  way1Tag_64 = _RAND_704[20:0];
  _RAND_705 = {1{`RANDOM}};
  way1Tag_65 = _RAND_705[20:0];
  _RAND_706 = {1{`RANDOM}};
  way1Tag_66 = _RAND_706[20:0];
  _RAND_707 = {1{`RANDOM}};
  way1Tag_67 = _RAND_707[20:0];
  _RAND_708 = {1{`RANDOM}};
  way1Tag_68 = _RAND_708[20:0];
  _RAND_709 = {1{`RANDOM}};
  way1Tag_69 = _RAND_709[20:0];
  _RAND_710 = {1{`RANDOM}};
  way1Tag_70 = _RAND_710[20:0];
  _RAND_711 = {1{`RANDOM}};
  way1Tag_71 = _RAND_711[20:0];
  _RAND_712 = {1{`RANDOM}};
  way1Tag_72 = _RAND_712[20:0];
  _RAND_713 = {1{`RANDOM}};
  way1Tag_73 = _RAND_713[20:0];
  _RAND_714 = {1{`RANDOM}};
  way1Tag_74 = _RAND_714[20:0];
  _RAND_715 = {1{`RANDOM}};
  way1Tag_75 = _RAND_715[20:0];
  _RAND_716 = {1{`RANDOM}};
  way1Tag_76 = _RAND_716[20:0];
  _RAND_717 = {1{`RANDOM}};
  way1Tag_77 = _RAND_717[20:0];
  _RAND_718 = {1{`RANDOM}};
  way1Tag_78 = _RAND_718[20:0];
  _RAND_719 = {1{`RANDOM}};
  way1Tag_79 = _RAND_719[20:0];
  _RAND_720 = {1{`RANDOM}};
  way1Tag_80 = _RAND_720[20:0];
  _RAND_721 = {1{`RANDOM}};
  way1Tag_81 = _RAND_721[20:0];
  _RAND_722 = {1{`RANDOM}};
  way1Tag_82 = _RAND_722[20:0];
  _RAND_723 = {1{`RANDOM}};
  way1Tag_83 = _RAND_723[20:0];
  _RAND_724 = {1{`RANDOM}};
  way1Tag_84 = _RAND_724[20:0];
  _RAND_725 = {1{`RANDOM}};
  way1Tag_85 = _RAND_725[20:0];
  _RAND_726 = {1{`RANDOM}};
  way1Tag_86 = _RAND_726[20:0];
  _RAND_727 = {1{`RANDOM}};
  way1Tag_87 = _RAND_727[20:0];
  _RAND_728 = {1{`RANDOM}};
  way1Tag_88 = _RAND_728[20:0];
  _RAND_729 = {1{`RANDOM}};
  way1Tag_89 = _RAND_729[20:0];
  _RAND_730 = {1{`RANDOM}};
  way1Tag_90 = _RAND_730[20:0];
  _RAND_731 = {1{`RANDOM}};
  way1Tag_91 = _RAND_731[20:0];
  _RAND_732 = {1{`RANDOM}};
  way1Tag_92 = _RAND_732[20:0];
  _RAND_733 = {1{`RANDOM}};
  way1Tag_93 = _RAND_733[20:0];
  _RAND_734 = {1{`RANDOM}};
  way1Tag_94 = _RAND_734[20:0];
  _RAND_735 = {1{`RANDOM}};
  way1Tag_95 = _RAND_735[20:0];
  _RAND_736 = {1{`RANDOM}};
  way1Tag_96 = _RAND_736[20:0];
  _RAND_737 = {1{`RANDOM}};
  way1Tag_97 = _RAND_737[20:0];
  _RAND_738 = {1{`RANDOM}};
  way1Tag_98 = _RAND_738[20:0];
  _RAND_739 = {1{`RANDOM}};
  way1Tag_99 = _RAND_739[20:0];
  _RAND_740 = {1{`RANDOM}};
  way1Tag_100 = _RAND_740[20:0];
  _RAND_741 = {1{`RANDOM}};
  way1Tag_101 = _RAND_741[20:0];
  _RAND_742 = {1{`RANDOM}};
  way1Tag_102 = _RAND_742[20:0];
  _RAND_743 = {1{`RANDOM}};
  way1Tag_103 = _RAND_743[20:0];
  _RAND_744 = {1{`RANDOM}};
  way1Tag_104 = _RAND_744[20:0];
  _RAND_745 = {1{`RANDOM}};
  way1Tag_105 = _RAND_745[20:0];
  _RAND_746 = {1{`RANDOM}};
  way1Tag_106 = _RAND_746[20:0];
  _RAND_747 = {1{`RANDOM}};
  way1Tag_107 = _RAND_747[20:0];
  _RAND_748 = {1{`RANDOM}};
  way1Tag_108 = _RAND_748[20:0];
  _RAND_749 = {1{`RANDOM}};
  way1Tag_109 = _RAND_749[20:0];
  _RAND_750 = {1{`RANDOM}};
  way1Tag_110 = _RAND_750[20:0];
  _RAND_751 = {1{`RANDOM}};
  way1Tag_111 = _RAND_751[20:0];
  _RAND_752 = {1{`RANDOM}};
  way1Tag_112 = _RAND_752[20:0];
  _RAND_753 = {1{`RANDOM}};
  way1Tag_113 = _RAND_753[20:0];
  _RAND_754 = {1{`RANDOM}};
  way1Tag_114 = _RAND_754[20:0];
  _RAND_755 = {1{`RANDOM}};
  way1Tag_115 = _RAND_755[20:0];
  _RAND_756 = {1{`RANDOM}};
  way1Tag_116 = _RAND_756[20:0];
  _RAND_757 = {1{`RANDOM}};
  way1Tag_117 = _RAND_757[20:0];
  _RAND_758 = {1{`RANDOM}};
  way1Tag_118 = _RAND_758[20:0];
  _RAND_759 = {1{`RANDOM}};
  way1Tag_119 = _RAND_759[20:0];
  _RAND_760 = {1{`RANDOM}};
  way1Tag_120 = _RAND_760[20:0];
  _RAND_761 = {1{`RANDOM}};
  way1Tag_121 = _RAND_761[20:0];
  _RAND_762 = {1{`RANDOM}};
  way1Tag_122 = _RAND_762[20:0];
  _RAND_763 = {1{`RANDOM}};
  way1Tag_123 = _RAND_763[20:0];
  _RAND_764 = {1{`RANDOM}};
  way1Tag_124 = _RAND_764[20:0];
  _RAND_765 = {1{`RANDOM}};
  way1Tag_125 = _RAND_765[20:0];
  _RAND_766 = {1{`RANDOM}};
  way1Tag_126 = _RAND_766[20:0];
  _RAND_767 = {1{`RANDOM}};
  way1Tag_127 = _RAND_767[20:0];
  _RAND_768 = {1{`RANDOM}};
  way1Age_0 = _RAND_768[0:0];
  _RAND_769 = {1{`RANDOM}};
  way1Age_1 = _RAND_769[0:0];
  _RAND_770 = {1{`RANDOM}};
  way1Age_2 = _RAND_770[0:0];
  _RAND_771 = {1{`RANDOM}};
  way1Age_3 = _RAND_771[0:0];
  _RAND_772 = {1{`RANDOM}};
  way1Age_4 = _RAND_772[0:0];
  _RAND_773 = {1{`RANDOM}};
  way1Age_5 = _RAND_773[0:0];
  _RAND_774 = {1{`RANDOM}};
  way1Age_6 = _RAND_774[0:0];
  _RAND_775 = {1{`RANDOM}};
  way1Age_7 = _RAND_775[0:0];
  _RAND_776 = {1{`RANDOM}};
  way1Age_8 = _RAND_776[0:0];
  _RAND_777 = {1{`RANDOM}};
  way1Age_9 = _RAND_777[0:0];
  _RAND_778 = {1{`RANDOM}};
  way1Age_10 = _RAND_778[0:0];
  _RAND_779 = {1{`RANDOM}};
  way1Age_11 = _RAND_779[0:0];
  _RAND_780 = {1{`RANDOM}};
  way1Age_12 = _RAND_780[0:0];
  _RAND_781 = {1{`RANDOM}};
  way1Age_13 = _RAND_781[0:0];
  _RAND_782 = {1{`RANDOM}};
  way1Age_14 = _RAND_782[0:0];
  _RAND_783 = {1{`RANDOM}};
  way1Age_15 = _RAND_783[0:0];
  _RAND_784 = {1{`RANDOM}};
  way1Age_16 = _RAND_784[0:0];
  _RAND_785 = {1{`RANDOM}};
  way1Age_17 = _RAND_785[0:0];
  _RAND_786 = {1{`RANDOM}};
  way1Age_18 = _RAND_786[0:0];
  _RAND_787 = {1{`RANDOM}};
  way1Age_19 = _RAND_787[0:0];
  _RAND_788 = {1{`RANDOM}};
  way1Age_20 = _RAND_788[0:0];
  _RAND_789 = {1{`RANDOM}};
  way1Age_21 = _RAND_789[0:0];
  _RAND_790 = {1{`RANDOM}};
  way1Age_22 = _RAND_790[0:0];
  _RAND_791 = {1{`RANDOM}};
  way1Age_23 = _RAND_791[0:0];
  _RAND_792 = {1{`RANDOM}};
  way1Age_24 = _RAND_792[0:0];
  _RAND_793 = {1{`RANDOM}};
  way1Age_25 = _RAND_793[0:0];
  _RAND_794 = {1{`RANDOM}};
  way1Age_26 = _RAND_794[0:0];
  _RAND_795 = {1{`RANDOM}};
  way1Age_27 = _RAND_795[0:0];
  _RAND_796 = {1{`RANDOM}};
  way1Age_28 = _RAND_796[0:0];
  _RAND_797 = {1{`RANDOM}};
  way1Age_29 = _RAND_797[0:0];
  _RAND_798 = {1{`RANDOM}};
  way1Age_30 = _RAND_798[0:0];
  _RAND_799 = {1{`RANDOM}};
  way1Age_31 = _RAND_799[0:0];
  _RAND_800 = {1{`RANDOM}};
  way1Age_32 = _RAND_800[0:0];
  _RAND_801 = {1{`RANDOM}};
  way1Age_33 = _RAND_801[0:0];
  _RAND_802 = {1{`RANDOM}};
  way1Age_34 = _RAND_802[0:0];
  _RAND_803 = {1{`RANDOM}};
  way1Age_35 = _RAND_803[0:0];
  _RAND_804 = {1{`RANDOM}};
  way1Age_36 = _RAND_804[0:0];
  _RAND_805 = {1{`RANDOM}};
  way1Age_37 = _RAND_805[0:0];
  _RAND_806 = {1{`RANDOM}};
  way1Age_38 = _RAND_806[0:0];
  _RAND_807 = {1{`RANDOM}};
  way1Age_39 = _RAND_807[0:0];
  _RAND_808 = {1{`RANDOM}};
  way1Age_40 = _RAND_808[0:0];
  _RAND_809 = {1{`RANDOM}};
  way1Age_41 = _RAND_809[0:0];
  _RAND_810 = {1{`RANDOM}};
  way1Age_42 = _RAND_810[0:0];
  _RAND_811 = {1{`RANDOM}};
  way1Age_43 = _RAND_811[0:0];
  _RAND_812 = {1{`RANDOM}};
  way1Age_44 = _RAND_812[0:0];
  _RAND_813 = {1{`RANDOM}};
  way1Age_45 = _RAND_813[0:0];
  _RAND_814 = {1{`RANDOM}};
  way1Age_46 = _RAND_814[0:0];
  _RAND_815 = {1{`RANDOM}};
  way1Age_47 = _RAND_815[0:0];
  _RAND_816 = {1{`RANDOM}};
  way1Age_48 = _RAND_816[0:0];
  _RAND_817 = {1{`RANDOM}};
  way1Age_49 = _RAND_817[0:0];
  _RAND_818 = {1{`RANDOM}};
  way1Age_50 = _RAND_818[0:0];
  _RAND_819 = {1{`RANDOM}};
  way1Age_51 = _RAND_819[0:0];
  _RAND_820 = {1{`RANDOM}};
  way1Age_52 = _RAND_820[0:0];
  _RAND_821 = {1{`RANDOM}};
  way1Age_53 = _RAND_821[0:0];
  _RAND_822 = {1{`RANDOM}};
  way1Age_54 = _RAND_822[0:0];
  _RAND_823 = {1{`RANDOM}};
  way1Age_55 = _RAND_823[0:0];
  _RAND_824 = {1{`RANDOM}};
  way1Age_56 = _RAND_824[0:0];
  _RAND_825 = {1{`RANDOM}};
  way1Age_57 = _RAND_825[0:0];
  _RAND_826 = {1{`RANDOM}};
  way1Age_58 = _RAND_826[0:0];
  _RAND_827 = {1{`RANDOM}};
  way1Age_59 = _RAND_827[0:0];
  _RAND_828 = {1{`RANDOM}};
  way1Age_60 = _RAND_828[0:0];
  _RAND_829 = {1{`RANDOM}};
  way1Age_61 = _RAND_829[0:0];
  _RAND_830 = {1{`RANDOM}};
  way1Age_62 = _RAND_830[0:0];
  _RAND_831 = {1{`RANDOM}};
  way1Age_63 = _RAND_831[0:0];
  _RAND_832 = {1{`RANDOM}};
  way1Age_64 = _RAND_832[0:0];
  _RAND_833 = {1{`RANDOM}};
  way1Age_65 = _RAND_833[0:0];
  _RAND_834 = {1{`RANDOM}};
  way1Age_66 = _RAND_834[0:0];
  _RAND_835 = {1{`RANDOM}};
  way1Age_67 = _RAND_835[0:0];
  _RAND_836 = {1{`RANDOM}};
  way1Age_68 = _RAND_836[0:0];
  _RAND_837 = {1{`RANDOM}};
  way1Age_69 = _RAND_837[0:0];
  _RAND_838 = {1{`RANDOM}};
  way1Age_70 = _RAND_838[0:0];
  _RAND_839 = {1{`RANDOM}};
  way1Age_71 = _RAND_839[0:0];
  _RAND_840 = {1{`RANDOM}};
  way1Age_72 = _RAND_840[0:0];
  _RAND_841 = {1{`RANDOM}};
  way1Age_73 = _RAND_841[0:0];
  _RAND_842 = {1{`RANDOM}};
  way1Age_74 = _RAND_842[0:0];
  _RAND_843 = {1{`RANDOM}};
  way1Age_75 = _RAND_843[0:0];
  _RAND_844 = {1{`RANDOM}};
  way1Age_76 = _RAND_844[0:0];
  _RAND_845 = {1{`RANDOM}};
  way1Age_77 = _RAND_845[0:0];
  _RAND_846 = {1{`RANDOM}};
  way1Age_78 = _RAND_846[0:0];
  _RAND_847 = {1{`RANDOM}};
  way1Age_79 = _RAND_847[0:0];
  _RAND_848 = {1{`RANDOM}};
  way1Age_80 = _RAND_848[0:0];
  _RAND_849 = {1{`RANDOM}};
  way1Age_81 = _RAND_849[0:0];
  _RAND_850 = {1{`RANDOM}};
  way1Age_82 = _RAND_850[0:0];
  _RAND_851 = {1{`RANDOM}};
  way1Age_83 = _RAND_851[0:0];
  _RAND_852 = {1{`RANDOM}};
  way1Age_84 = _RAND_852[0:0];
  _RAND_853 = {1{`RANDOM}};
  way1Age_85 = _RAND_853[0:0];
  _RAND_854 = {1{`RANDOM}};
  way1Age_86 = _RAND_854[0:0];
  _RAND_855 = {1{`RANDOM}};
  way1Age_87 = _RAND_855[0:0];
  _RAND_856 = {1{`RANDOM}};
  way1Age_88 = _RAND_856[0:0];
  _RAND_857 = {1{`RANDOM}};
  way1Age_89 = _RAND_857[0:0];
  _RAND_858 = {1{`RANDOM}};
  way1Age_90 = _RAND_858[0:0];
  _RAND_859 = {1{`RANDOM}};
  way1Age_91 = _RAND_859[0:0];
  _RAND_860 = {1{`RANDOM}};
  way1Age_92 = _RAND_860[0:0];
  _RAND_861 = {1{`RANDOM}};
  way1Age_93 = _RAND_861[0:0];
  _RAND_862 = {1{`RANDOM}};
  way1Age_94 = _RAND_862[0:0];
  _RAND_863 = {1{`RANDOM}};
  way1Age_95 = _RAND_863[0:0];
  _RAND_864 = {1{`RANDOM}};
  way1Age_96 = _RAND_864[0:0];
  _RAND_865 = {1{`RANDOM}};
  way1Age_97 = _RAND_865[0:0];
  _RAND_866 = {1{`RANDOM}};
  way1Age_98 = _RAND_866[0:0];
  _RAND_867 = {1{`RANDOM}};
  way1Age_99 = _RAND_867[0:0];
  _RAND_868 = {1{`RANDOM}};
  way1Age_100 = _RAND_868[0:0];
  _RAND_869 = {1{`RANDOM}};
  way1Age_101 = _RAND_869[0:0];
  _RAND_870 = {1{`RANDOM}};
  way1Age_102 = _RAND_870[0:0];
  _RAND_871 = {1{`RANDOM}};
  way1Age_103 = _RAND_871[0:0];
  _RAND_872 = {1{`RANDOM}};
  way1Age_104 = _RAND_872[0:0];
  _RAND_873 = {1{`RANDOM}};
  way1Age_105 = _RAND_873[0:0];
  _RAND_874 = {1{`RANDOM}};
  way1Age_106 = _RAND_874[0:0];
  _RAND_875 = {1{`RANDOM}};
  way1Age_107 = _RAND_875[0:0];
  _RAND_876 = {1{`RANDOM}};
  way1Age_108 = _RAND_876[0:0];
  _RAND_877 = {1{`RANDOM}};
  way1Age_109 = _RAND_877[0:0];
  _RAND_878 = {1{`RANDOM}};
  way1Age_110 = _RAND_878[0:0];
  _RAND_879 = {1{`RANDOM}};
  way1Age_111 = _RAND_879[0:0];
  _RAND_880 = {1{`RANDOM}};
  way1Age_112 = _RAND_880[0:0];
  _RAND_881 = {1{`RANDOM}};
  way1Age_113 = _RAND_881[0:0];
  _RAND_882 = {1{`RANDOM}};
  way1Age_114 = _RAND_882[0:0];
  _RAND_883 = {1{`RANDOM}};
  way1Age_115 = _RAND_883[0:0];
  _RAND_884 = {1{`RANDOM}};
  way1Age_116 = _RAND_884[0:0];
  _RAND_885 = {1{`RANDOM}};
  way1Age_117 = _RAND_885[0:0];
  _RAND_886 = {1{`RANDOM}};
  way1Age_118 = _RAND_886[0:0];
  _RAND_887 = {1{`RANDOM}};
  way1Age_119 = _RAND_887[0:0];
  _RAND_888 = {1{`RANDOM}};
  way1Age_120 = _RAND_888[0:0];
  _RAND_889 = {1{`RANDOM}};
  way1Age_121 = _RAND_889[0:0];
  _RAND_890 = {1{`RANDOM}};
  way1Age_122 = _RAND_890[0:0];
  _RAND_891 = {1{`RANDOM}};
  way1Age_123 = _RAND_891[0:0];
  _RAND_892 = {1{`RANDOM}};
  way1Age_124 = _RAND_892[0:0];
  _RAND_893 = {1{`RANDOM}};
  way1Age_125 = _RAND_893[0:0];
  _RAND_894 = {1{`RANDOM}};
  way1Age_126 = _RAND_894[0:0];
  _RAND_895 = {1{`RANDOM}};
  way1Age_127 = _RAND_895[0:0];
  _RAND_896 = {1{`RANDOM}};
  way1Dirty_0 = _RAND_896[0:0];
  _RAND_897 = {1{`RANDOM}};
  way1Dirty_1 = _RAND_897[0:0];
  _RAND_898 = {1{`RANDOM}};
  way1Dirty_2 = _RAND_898[0:0];
  _RAND_899 = {1{`RANDOM}};
  way1Dirty_3 = _RAND_899[0:0];
  _RAND_900 = {1{`RANDOM}};
  way1Dirty_4 = _RAND_900[0:0];
  _RAND_901 = {1{`RANDOM}};
  way1Dirty_5 = _RAND_901[0:0];
  _RAND_902 = {1{`RANDOM}};
  way1Dirty_6 = _RAND_902[0:0];
  _RAND_903 = {1{`RANDOM}};
  way1Dirty_7 = _RAND_903[0:0];
  _RAND_904 = {1{`RANDOM}};
  way1Dirty_8 = _RAND_904[0:0];
  _RAND_905 = {1{`RANDOM}};
  way1Dirty_9 = _RAND_905[0:0];
  _RAND_906 = {1{`RANDOM}};
  way1Dirty_10 = _RAND_906[0:0];
  _RAND_907 = {1{`RANDOM}};
  way1Dirty_11 = _RAND_907[0:0];
  _RAND_908 = {1{`RANDOM}};
  way1Dirty_12 = _RAND_908[0:0];
  _RAND_909 = {1{`RANDOM}};
  way1Dirty_13 = _RAND_909[0:0];
  _RAND_910 = {1{`RANDOM}};
  way1Dirty_14 = _RAND_910[0:0];
  _RAND_911 = {1{`RANDOM}};
  way1Dirty_15 = _RAND_911[0:0];
  _RAND_912 = {1{`RANDOM}};
  way1Dirty_16 = _RAND_912[0:0];
  _RAND_913 = {1{`RANDOM}};
  way1Dirty_17 = _RAND_913[0:0];
  _RAND_914 = {1{`RANDOM}};
  way1Dirty_18 = _RAND_914[0:0];
  _RAND_915 = {1{`RANDOM}};
  way1Dirty_19 = _RAND_915[0:0];
  _RAND_916 = {1{`RANDOM}};
  way1Dirty_20 = _RAND_916[0:0];
  _RAND_917 = {1{`RANDOM}};
  way1Dirty_21 = _RAND_917[0:0];
  _RAND_918 = {1{`RANDOM}};
  way1Dirty_22 = _RAND_918[0:0];
  _RAND_919 = {1{`RANDOM}};
  way1Dirty_23 = _RAND_919[0:0];
  _RAND_920 = {1{`RANDOM}};
  way1Dirty_24 = _RAND_920[0:0];
  _RAND_921 = {1{`RANDOM}};
  way1Dirty_25 = _RAND_921[0:0];
  _RAND_922 = {1{`RANDOM}};
  way1Dirty_26 = _RAND_922[0:0];
  _RAND_923 = {1{`RANDOM}};
  way1Dirty_27 = _RAND_923[0:0];
  _RAND_924 = {1{`RANDOM}};
  way1Dirty_28 = _RAND_924[0:0];
  _RAND_925 = {1{`RANDOM}};
  way1Dirty_29 = _RAND_925[0:0];
  _RAND_926 = {1{`RANDOM}};
  way1Dirty_30 = _RAND_926[0:0];
  _RAND_927 = {1{`RANDOM}};
  way1Dirty_31 = _RAND_927[0:0];
  _RAND_928 = {1{`RANDOM}};
  way1Dirty_32 = _RAND_928[0:0];
  _RAND_929 = {1{`RANDOM}};
  way1Dirty_33 = _RAND_929[0:0];
  _RAND_930 = {1{`RANDOM}};
  way1Dirty_34 = _RAND_930[0:0];
  _RAND_931 = {1{`RANDOM}};
  way1Dirty_35 = _RAND_931[0:0];
  _RAND_932 = {1{`RANDOM}};
  way1Dirty_36 = _RAND_932[0:0];
  _RAND_933 = {1{`RANDOM}};
  way1Dirty_37 = _RAND_933[0:0];
  _RAND_934 = {1{`RANDOM}};
  way1Dirty_38 = _RAND_934[0:0];
  _RAND_935 = {1{`RANDOM}};
  way1Dirty_39 = _RAND_935[0:0];
  _RAND_936 = {1{`RANDOM}};
  way1Dirty_40 = _RAND_936[0:0];
  _RAND_937 = {1{`RANDOM}};
  way1Dirty_41 = _RAND_937[0:0];
  _RAND_938 = {1{`RANDOM}};
  way1Dirty_42 = _RAND_938[0:0];
  _RAND_939 = {1{`RANDOM}};
  way1Dirty_43 = _RAND_939[0:0];
  _RAND_940 = {1{`RANDOM}};
  way1Dirty_44 = _RAND_940[0:0];
  _RAND_941 = {1{`RANDOM}};
  way1Dirty_45 = _RAND_941[0:0];
  _RAND_942 = {1{`RANDOM}};
  way1Dirty_46 = _RAND_942[0:0];
  _RAND_943 = {1{`RANDOM}};
  way1Dirty_47 = _RAND_943[0:0];
  _RAND_944 = {1{`RANDOM}};
  way1Dirty_48 = _RAND_944[0:0];
  _RAND_945 = {1{`RANDOM}};
  way1Dirty_49 = _RAND_945[0:0];
  _RAND_946 = {1{`RANDOM}};
  way1Dirty_50 = _RAND_946[0:0];
  _RAND_947 = {1{`RANDOM}};
  way1Dirty_51 = _RAND_947[0:0];
  _RAND_948 = {1{`RANDOM}};
  way1Dirty_52 = _RAND_948[0:0];
  _RAND_949 = {1{`RANDOM}};
  way1Dirty_53 = _RAND_949[0:0];
  _RAND_950 = {1{`RANDOM}};
  way1Dirty_54 = _RAND_950[0:0];
  _RAND_951 = {1{`RANDOM}};
  way1Dirty_55 = _RAND_951[0:0];
  _RAND_952 = {1{`RANDOM}};
  way1Dirty_56 = _RAND_952[0:0];
  _RAND_953 = {1{`RANDOM}};
  way1Dirty_57 = _RAND_953[0:0];
  _RAND_954 = {1{`RANDOM}};
  way1Dirty_58 = _RAND_954[0:0];
  _RAND_955 = {1{`RANDOM}};
  way1Dirty_59 = _RAND_955[0:0];
  _RAND_956 = {1{`RANDOM}};
  way1Dirty_60 = _RAND_956[0:0];
  _RAND_957 = {1{`RANDOM}};
  way1Dirty_61 = _RAND_957[0:0];
  _RAND_958 = {1{`RANDOM}};
  way1Dirty_62 = _RAND_958[0:0];
  _RAND_959 = {1{`RANDOM}};
  way1Dirty_63 = _RAND_959[0:0];
  _RAND_960 = {1{`RANDOM}};
  way1Dirty_64 = _RAND_960[0:0];
  _RAND_961 = {1{`RANDOM}};
  way1Dirty_65 = _RAND_961[0:0];
  _RAND_962 = {1{`RANDOM}};
  way1Dirty_66 = _RAND_962[0:0];
  _RAND_963 = {1{`RANDOM}};
  way1Dirty_67 = _RAND_963[0:0];
  _RAND_964 = {1{`RANDOM}};
  way1Dirty_68 = _RAND_964[0:0];
  _RAND_965 = {1{`RANDOM}};
  way1Dirty_69 = _RAND_965[0:0];
  _RAND_966 = {1{`RANDOM}};
  way1Dirty_70 = _RAND_966[0:0];
  _RAND_967 = {1{`RANDOM}};
  way1Dirty_71 = _RAND_967[0:0];
  _RAND_968 = {1{`RANDOM}};
  way1Dirty_72 = _RAND_968[0:0];
  _RAND_969 = {1{`RANDOM}};
  way1Dirty_73 = _RAND_969[0:0];
  _RAND_970 = {1{`RANDOM}};
  way1Dirty_74 = _RAND_970[0:0];
  _RAND_971 = {1{`RANDOM}};
  way1Dirty_75 = _RAND_971[0:0];
  _RAND_972 = {1{`RANDOM}};
  way1Dirty_76 = _RAND_972[0:0];
  _RAND_973 = {1{`RANDOM}};
  way1Dirty_77 = _RAND_973[0:0];
  _RAND_974 = {1{`RANDOM}};
  way1Dirty_78 = _RAND_974[0:0];
  _RAND_975 = {1{`RANDOM}};
  way1Dirty_79 = _RAND_975[0:0];
  _RAND_976 = {1{`RANDOM}};
  way1Dirty_80 = _RAND_976[0:0];
  _RAND_977 = {1{`RANDOM}};
  way1Dirty_81 = _RAND_977[0:0];
  _RAND_978 = {1{`RANDOM}};
  way1Dirty_82 = _RAND_978[0:0];
  _RAND_979 = {1{`RANDOM}};
  way1Dirty_83 = _RAND_979[0:0];
  _RAND_980 = {1{`RANDOM}};
  way1Dirty_84 = _RAND_980[0:0];
  _RAND_981 = {1{`RANDOM}};
  way1Dirty_85 = _RAND_981[0:0];
  _RAND_982 = {1{`RANDOM}};
  way1Dirty_86 = _RAND_982[0:0];
  _RAND_983 = {1{`RANDOM}};
  way1Dirty_87 = _RAND_983[0:0];
  _RAND_984 = {1{`RANDOM}};
  way1Dirty_88 = _RAND_984[0:0];
  _RAND_985 = {1{`RANDOM}};
  way1Dirty_89 = _RAND_985[0:0];
  _RAND_986 = {1{`RANDOM}};
  way1Dirty_90 = _RAND_986[0:0];
  _RAND_987 = {1{`RANDOM}};
  way1Dirty_91 = _RAND_987[0:0];
  _RAND_988 = {1{`RANDOM}};
  way1Dirty_92 = _RAND_988[0:0];
  _RAND_989 = {1{`RANDOM}};
  way1Dirty_93 = _RAND_989[0:0];
  _RAND_990 = {1{`RANDOM}};
  way1Dirty_94 = _RAND_990[0:0];
  _RAND_991 = {1{`RANDOM}};
  way1Dirty_95 = _RAND_991[0:0];
  _RAND_992 = {1{`RANDOM}};
  way1Dirty_96 = _RAND_992[0:0];
  _RAND_993 = {1{`RANDOM}};
  way1Dirty_97 = _RAND_993[0:0];
  _RAND_994 = {1{`RANDOM}};
  way1Dirty_98 = _RAND_994[0:0];
  _RAND_995 = {1{`RANDOM}};
  way1Dirty_99 = _RAND_995[0:0];
  _RAND_996 = {1{`RANDOM}};
  way1Dirty_100 = _RAND_996[0:0];
  _RAND_997 = {1{`RANDOM}};
  way1Dirty_101 = _RAND_997[0:0];
  _RAND_998 = {1{`RANDOM}};
  way1Dirty_102 = _RAND_998[0:0];
  _RAND_999 = {1{`RANDOM}};
  way1Dirty_103 = _RAND_999[0:0];
  _RAND_1000 = {1{`RANDOM}};
  way1Dirty_104 = _RAND_1000[0:0];
  _RAND_1001 = {1{`RANDOM}};
  way1Dirty_105 = _RAND_1001[0:0];
  _RAND_1002 = {1{`RANDOM}};
  way1Dirty_106 = _RAND_1002[0:0];
  _RAND_1003 = {1{`RANDOM}};
  way1Dirty_107 = _RAND_1003[0:0];
  _RAND_1004 = {1{`RANDOM}};
  way1Dirty_108 = _RAND_1004[0:0];
  _RAND_1005 = {1{`RANDOM}};
  way1Dirty_109 = _RAND_1005[0:0];
  _RAND_1006 = {1{`RANDOM}};
  way1Dirty_110 = _RAND_1006[0:0];
  _RAND_1007 = {1{`RANDOM}};
  way1Dirty_111 = _RAND_1007[0:0];
  _RAND_1008 = {1{`RANDOM}};
  way1Dirty_112 = _RAND_1008[0:0];
  _RAND_1009 = {1{`RANDOM}};
  way1Dirty_113 = _RAND_1009[0:0];
  _RAND_1010 = {1{`RANDOM}};
  way1Dirty_114 = _RAND_1010[0:0];
  _RAND_1011 = {1{`RANDOM}};
  way1Dirty_115 = _RAND_1011[0:0];
  _RAND_1012 = {1{`RANDOM}};
  way1Dirty_116 = _RAND_1012[0:0];
  _RAND_1013 = {1{`RANDOM}};
  way1Dirty_117 = _RAND_1013[0:0];
  _RAND_1014 = {1{`RANDOM}};
  way1Dirty_118 = _RAND_1014[0:0];
  _RAND_1015 = {1{`RANDOM}};
  way1Dirty_119 = _RAND_1015[0:0];
  _RAND_1016 = {1{`RANDOM}};
  way1Dirty_120 = _RAND_1016[0:0];
  _RAND_1017 = {1{`RANDOM}};
  way1Dirty_121 = _RAND_1017[0:0];
  _RAND_1018 = {1{`RANDOM}};
  way1Dirty_122 = _RAND_1018[0:0];
  _RAND_1019 = {1{`RANDOM}};
  way1Dirty_123 = _RAND_1019[0:0];
  _RAND_1020 = {1{`RANDOM}};
  way1Dirty_124 = _RAND_1020[0:0];
  _RAND_1021 = {1{`RANDOM}};
  way1Dirty_125 = _RAND_1021[0:0];
  _RAND_1022 = {1{`RANDOM}};
  way1Dirty_126 = _RAND_1022[0:0];
  _RAND_1023 = {1{`RANDOM}};
  way1Dirty_127 = _RAND_1023[0:0];
  _RAND_1024 = {1{`RANDOM}};
  state = _RAND_1024[2:0];
  _RAND_1025 = {1{`RANDOM}};
  hitEn = _RAND_1025[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AxiLite2Axi(
  input          clock,
  input          reset,
  input          io_out_aw_ready,
  output         io_out_aw_valid,
  output [31:0]  io_out_aw_bits_addr,
  input          io_out_w_ready,
  output         io_out_w_valid,
  output [63:0]  io_out_w_bits_data,
  output [7:0]   io_out_w_bits_strb,
  output         io_out_w_bits_last,
  output         io_out_b_ready,
  input          io_out_b_valid,
  input          io_out_ar_ready,
  output         io_out_ar_valid,
  output [31:0]  io_out_ar_bits_addr,
  output         io_out_r_ready,
  input          io_out_r_valid,
  input  [63:0]  io_out_r_bits_data,
  input          io_out_r_bits_last,
  input          io_imem_inst_valid,
  output         io_imem_inst_ready,
  input  [31:0]  io_imem_inst_addr,
  output [127:0] io_imem_inst_read,
  input          io_dmem_data_valid,
  output         io_dmem_data_ready,
  input          io_dmem_data_req,
  input  [31:0]  io_dmem_data_addr,
  input  [7:0]   io_dmem_data_strb,
  output [127:0] io_dmem_data_read,
  input  [127:0] io_dmem_data_write
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  wire  data_ren = io_dmem_data_valid & ~io_dmem_data_req; // @[Axi.scala 29:30]
  wire  data_wen = io_dmem_data_valid & io_dmem_data_req; // @[Axi.scala 30:30]
  wire  ar_hs = io_out_ar_ready & io_out_ar_valid; // @[Axi.scala 32:28]
  wire  r_hs = io_out_r_valid & io_out_r_ready; // @[Axi.scala 33:26]
  wire  aw_hs = io_out_aw_ready & io_out_aw_valid; // @[Axi.scala 34:28]
  wire  w_hs = io_out_w_ready & io_out_w_valid; // @[Axi.scala 35:26]
  wire  b_hs = io_out_b_valid & io_out_b_ready; // @[Axi.scala 36:26]
  wire  r_done = r_hs & io_out_r_bits_last; // @[Axi.scala 38:21]
  wire  w_done = b_hs & io_out_w_bits_last; // @[Axi.scala 39:21]
  reg [2:0] r_state; // @[Axi.scala 43:24]
  reg [2:0] w_state; // @[Axi.scala 44:24]
  wire [2:0] _GEN_3 = r_done ? 3'h3 : r_state; // @[Axi.scala 66:20 67:17 43:24]
  wire [2:0] _GEN_4 = data_ren ? 3'h4 : 3'h0; // @[Axi.scala 74:23 75:17 78:17]
  wire [2:0] _GEN_5 = ar_hs ? 3'h5 : r_state; // @[Axi.scala 82:20 83:17 43:24]
  wire [2:0] _GEN_6 = r_done ? 3'h6 : r_state; // @[Axi.scala 87:21 88:17 43:24]
  wire [2:0] _GEN_7 = 3'h6 == r_state ? 3'h0 : r_state; // @[Axi.scala 52:20 92:15 43:24]
  wire [2:0] _GEN_8 = 3'h5 == r_state ? _GEN_6 : _GEN_7; // @[Axi.scala 52:20]
  wire [2:0] _GEN_9 = 3'h4 == r_state ? _GEN_5 : _GEN_8; // @[Axi.scala 52:20]
  wire [2:0] _GEN_10 = 3'h3 == r_state ? _GEN_4 : _GEN_9; // @[Axi.scala 52:20]
  wire [2:0] _GEN_16 = w_hs ? 3'h3 : w_state; // @[Axi.scala 109:18 110:17 44:24]
  wire [2:0] _GEN_17 = w_done ? 3'h4 : w_state; // @[Axi.scala 114:20 115:17 44:24]
  wire [2:0] _GEN_18 = 3'h4 == w_state ? 3'h0 : w_state; // @[Axi.scala 119:15 97:20 44:24]
  wire [2:0] _GEN_19 = 3'h3 == w_state ? _GEN_17 : _GEN_18; // @[Axi.scala 97:20]
  reg  data_ok; // @[Axi.scala 123:24]
  wire  _T_12 = w_state == 3'h4; // @[Axi.scala 124:29]
  wire  _GEN_23 = ~data_wen ? 1'h0 : data_ok; // @[Axi.scala 127:25 128:13 123:24]
  wire  _GEN_24 = data_wen & w_state == 3'h4 | _GEN_23; // @[Axi.scala 124:46 125:13]
  wire  _axi_addr_T = r_state == 3'h1; // @[Axi.scala 131:30]
  wire [31:0] _axi_addr_T_1 = io_imem_inst_addr & 32'hfffffff0; // @[Axi.scala 131:63]
  wire  _axi_addr_T_2 = r_state == 3'h4; // @[Axi.scala 132:31]
  wire [31:0] _axi_addr_T_3 = io_dmem_data_addr & 32'hfffffff0; // @[Axi.scala 132:64]
  wire [31:0] _axi_addr_T_4 = r_state == 3'h4 ? _axi_addr_T_3 : 32'h0; // @[Axi.scala 132:22]
  wire [31:0] _axi_waddr_T_1 = {io_dmem_data_addr[31:4],4'h8}; // @[Cat.scala 31:58]
  reg [63:0] inst_read_h; // @[Axi.scala 184:28]
  reg [63:0] inst_read_l; // @[Axi.scala 185:28]
  reg [63:0] data_read_h; // @[Axi.scala 186:28]
  reg [63:0] data_read_l; // @[Axi.scala 187:28]
  assign io_out_aw_valid = w_state == 3'h1; // @[Axi.scala 160:34]
  assign io_out_aw_bits_addr = data_ok ? _axi_waddr_T_1 : _axi_addr_T_3; // @[Axi.scala 158:22]
  assign io_out_w_valid = w_state == 3'h2; // @[Axi.scala 173:34]
  assign io_out_w_bits_data = data_ok ? io_dmem_data_write[127:64] : io_dmem_data_write[63:0]; // @[Axi.scala 174:29]
  assign io_out_w_bits_strb = io_dmem_data_strb; // @[Axi.scala 175:23]
  assign io_out_w_bits_last = 1'h1; // @[Axi.scala 176:23]
  assign io_out_b_ready = 1'h1; // @[Axi.scala 178:23]
  assign io_out_ar_valid = _axi_addr_T | _axi_addr_T_2; // @[Axi.scala 142:44]
  assign io_out_ar_bits_addr = r_state == 3'h1 ? _axi_addr_T_1 : _axi_addr_T_4; // @[Axi.scala 131:21]
  assign io_out_r_ready = 1'h1; // @[Axi.scala 155:15]
  assign io_imem_inst_ready = r_state == 3'h3; // @[Axi.scala 181:30]
  assign io_imem_inst_read = {inst_read_h,inst_read_l}; // @[Cat.scala 31:58]
  assign io_dmem_data_ready = r_state == 3'h6 | _T_12 & data_ok; // @[Axi.scala 182:47]
  assign io_dmem_data_read = {data_read_h,data_read_l}; // @[Cat.scala 31:58]
  always @(posedge clock) begin
    if (reset) begin // @[Axi.scala 43:24]
      r_state <= 3'h0; // @[Axi.scala 43:24]
    end else if (3'h0 == r_state) begin // @[Axi.scala 52:20]
      if (io_imem_inst_valid) begin // @[Axi.scala 54:22]
        r_state <= 3'h1; // @[Axi.scala 55:17]
      end else if (data_ren) begin // @[Axi.scala 56:30]
        r_state <= 3'h4; // @[Axi.scala 57:17]
      end
    end else if (3'h1 == r_state) begin // @[Axi.scala 52:20]
      if (ar_hs) begin // @[Axi.scala 61:19]
        r_state <= 3'h2; // @[Axi.scala 62:17]
      end
    end else if (3'h2 == r_state) begin // @[Axi.scala 52:20]
      r_state <= _GEN_3;
    end else begin
      r_state <= _GEN_10;
    end
    if (reset) begin // @[Axi.scala 44:24]
      w_state <= 3'h0; // @[Axi.scala 44:24]
    end else if (3'h0 == w_state) begin // @[Axi.scala 97:20]
      if (data_wen) begin // @[Axi.scala 99:22]
        w_state <= 3'h1; // @[Axi.scala 100:17]
      end
    end else if (3'h1 == w_state) begin // @[Axi.scala 97:20]
      if (aw_hs) begin // @[Axi.scala 104:19]
        w_state <= 3'h2; // @[Axi.scala 105:17]
      end
    end else if (3'h2 == w_state) begin // @[Axi.scala 97:20]
      w_state <= _GEN_16;
    end else begin
      w_state <= _GEN_19;
    end
    if (reset) begin // @[Axi.scala 123:24]
      data_ok <= 1'h0; // @[Axi.scala 123:24]
    end else begin
      data_ok <= _GEN_24;
    end
    if (reset) begin // @[Axi.scala 184:28]
      inst_read_h <= 64'h0; // @[Axi.scala 184:28]
    end else if (r_hs) begin // @[Axi.scala 189:15]
      if (io_out_r_bits_last) begin // @[Axi.scala 190:28]
        inst_read_h <= io_out_r_bits_data; // @[Axi.scala 191:19]
      end
    end
    if (reset) begin // @[Axi.scala 185:28]
      inst_read_l <= 64'h0; // @[Axi.scala 185:28]
    end else if (r_hs) begin // @[Axi.scala 189:15]
      if (!(io_out_r_bits_last)) begin // @[Axi.scala 190:28]
        inst_read_l <= io_out_r_bits_data; // @[Axi.scala 195:19]
      end
    end
    if (reset) begin // @[Axi.scala 186:28]
      data_read_h <= 64'h0; // @[Axi.scala 186:28]
    end else if (r_hs) begin // @[Axi.scala 189:15]
      if (io_out_r_bits_last) begin // @[Axi.scala 190:28]
        data_read_h <= io_out_r_bits_data; // @[Axi.scala 192:19]
      end
    end
    if (reset) begin // @[Axi.scala 187:28]
      data_read_l <= 64'h0; // @[Axi.scala 187:28]
    end else if (r_hs) begin // @[Axi.scala 189:15]
      if (!(io_out_r_bits_last)) begin // @[Axi.scala 190:28]
        data_read_l <= io_out_r_bits_data; // @[Axi.scala 196:19]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r_state = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  w_state = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  data_ok = _RAND_2[0:0];
  _RAND_3 = {2{`RANDOM}};
  inst_read_h = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  inst_read_l = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  data_read_h = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  data_read_l = _RAND_6[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SimTop(
  input         clock,
  input         reset,
  input  [63:0] io_logCtrl_log_begin,
  input  [63:0] io_logCtrl_log_end,
  input  [63:0] io_logCtrl_log_level,
  input         io_perfInfo_clean,
  input         io_perfInfo_dump,
  output        io_uart_out_valid,
  output [7:0]  io_uart_out_ch,
  output        io_uart_in_valid,
  input  [7:0]  io_uart_in_ch,
  input         io_memAXI_0_aw_ready,
  output        io_memAXI_0_aw_valid,
  output [31:0] io_memAXI_0_aw_bits_addr,
  output [2:0]  io_memAXI_0_aw_bits_prot,
  output [3:0]  io_memAXI_0_aw_bits_id,
  output        io_memAXI_0_aw_bits_user,
  output [7:0]  io_memAXI_0_aw_bits_len,
  output [2:0]  io_memAXI_0_aw_bits_size,
  output [1:0]  io_memAXI_0_aw_bits_burst,
  output        io_memAXI_0_aw_bits_lock,
  output [3:0]  io_memAXI_0_aw_bits_cache,
  output [3:0]  io_memAXI_0_aw_bits_qos,
  input         io_memAXI_0_w_ready,
  output        io_memAXI_0_w_valid,
  output [63:0] io_memAXI_0_w_bits_data[3:0],
  output [7:0]  io_memAXI_0_w_bits_strb,
  output        io_memAXI_0_w_bits_last,
  output        io_memAXI_0_b_ready,
  input         io_memAXI_0_b_valid,
  input  [1:0]  io_memAXI_0_b_bits_resp,
  input  [3:0]  io_memAXI_0_b_bits_id,
  input         io_memAXI_0_b_bits_user,
  input         io_memAXI_0_ar_ready,
  output        io_memAXI_0_ar_valid,
  output [31:0] io_memAXI_0_ar_bits_addr,
  output [2:0]  io_memAXI_0_ar_bits_prot,
  output [3:0]  io_memAXI_0_ar_bits_id,
  output        io_memAXI_0_ar_bits_user,
  output [7:0]  io_memAXI_0_ar_bits_len,
  output [2:0]  io_memAXI_0_ar_bits_size,
  output [1:0]  io_memAXI_0_ar_bits_burst,
  output        io_memAXI_0_ar_bits_lock,
  output [3:0]  io_memAXI_0_ar_bits_cache,
  output [3:0]  io_memAXI_0_ar_bits_qos,
  output        io_memAXI_0_r_ready,
  input         io_memAXI_0_r_valid,
  input  [1:0]  io_memAXI_0_r_bits_resp,
  input  [63:0] io_memAXI_0_r_bits_data[3:0],
  input  [3:0]  io_memAXI_0_r_bits_id,
  input         io_memAXI_0_r_bits_user,
  input         io_memAXI_0_r_bits_last
);
  wire  core_clock; // @[SimTop.scala 18:20]
  wire  core_reset; // @[SimTop.scala 18:20]
  wire  core_io_imem_inst_valid; // @[SimTop.scala 18:20]
  wire  core_io_imem_inst_ready; // @[SimTop.scala 18:20]
  wire [31:0] core_io_imem_inst_addr; // @[SimTop.scala 18:20]
  wire [31:0] core_io_imem_inst_read; // @[SimTop.scala 18:20]
  wire  core_io_dmem_data_valid; // @[SimTop.scala 18:20]
  wire  core_io_dmem_data_ready; // @[SimTop.scala 18:20]
  wire  core_io_dmem_data_req; // @[SimTop.scala 18:20]
  wire [31:0] core_io_dmem_data_addr; // @[SimTop.scala 18:20]
  wire [1:0] core_io_dmem_data_size; // @[SimTop.scala 18:20]
  wire [7:0] core_io_dmem_data_strb; // @[SimTop.scala 18:20]
  wire [63:0] core_io_dmem_data_read; // @[SimTop.scala 18:20]
  wire [127:0] core_io_dmem_data_write; // @[SimTop.scala 18:20]
  wire  icache_clock; // @[SimTop.scala 19:22]
  wire  icache_reset; // @[SimTop.scala 19:22]
  wire  icache_io_imem_inst_valid; // @[SimTop.scala 19:22]
  wire  icache_io_imem_inst_ready; // @[SimTop.scala 19:22]
  wire [31:0] icache_io_imem_inst_addr; // @[SimTop.scala 19:22]
  wire [31:0] icache_io_imem_inst_read; // @[SimTop.scala 19:22]
  wire  icache_io_out_inst_valid; // @[SimTop.scala 19:22]
  wire  icache_io_out_inst_ready; // @[SimTop.scala 19:22]
  wire [31:0] icache_io_out_inst_addr; // @[SimTop.scala 19:22]
  wire [127:0] icache_io_out_inst_read; // @[SimTop.scala 19:22]
  wire  dcache_clock; // @[SimTop.scala 20:22]
  wire  dcache_reset; // @[SimTop.scala 20:22]
  wire  dcache_io_dmem_data_valid; // @[SimTop.scala 20:22]
  wire  dcache_io_dmem_data_ready; // @[SimTop.scala 20:22]
  wire  dcache_io_dmem_data_req; // @[SimTop.scala 20:22]
  wire [31:0] dcache_io_dmem_data_addr; // @[SimTop.scala 20:22]
  wire [1:0] dcache_io_dmem_data_size; // @[SimTop.scala 20:22]
  wire [7:0] dcache_io_dmem_data_strb; // @[SimTop.scala 20:22]
  wire [63:0] dcache_io_dmem_data_read; // @[SimTop.scala 20:22]
  wire [127:0] dcache_io_dmem_data_write; // @[SimTop.scala 20:22]
  wire  dcache_io_out_data_valid; // @[SimTop.scala 20:22]
  wire  dcache_io_out_data_ready; // @[SimTop.scala 20:22]
  wire  dcache_io_out_data_req; // @[SimTop.scala 20:22]
  wire [31:0] dcache_io_out_data_addr; // @[SimTop.scala 20:22]
  wire [7:0] dcache_io_out_data_strb; // @[SimTop.scala 20:22]
  wire [127:0] dcache_io_out_data_read; // @[SimTop.scala 20:22]
  wire [127:0] dcache_io_out_data_write; // @[SimTop.scala 20:22]
  wire  top_clock; // @[SimTop.scala 23:19]
  wire  top_reset; // @[SimTop.scala 23:19]
  wire  top_io_out_aw_ready; // @[SimTop.scala 23:19]
  wire  top_io_out_aw_valid; // @[SimTop.scala 23:19]
  wire [31:0] top_io_out_aw_bits_addr; // @[SimTop.scala 23:19]
  wire  top_io_out_w_ready; // @[SimTop.scala 23:19]
  wire  top_io_out_w_valid; // @[SimTop.scala 23:19]
  wire [63:0] top_io_out_w_bits_data; // @[SimTop.scala 23:19]
  wire [7:0] top_io_out_w_bits_strb; // @[SimTop.scala 23:19]
  wire  top_io_out_w_bits_last; // @[SimTop.scala 23:19]
  wire  top_io_out_b_ready; // @[SimTop.scala 23:19]
  wire  top_io_out_b_valid; // @[SimTop.scala 23:19]
  wire  top_io_out_ar_ready; // @[SimTop.scala 23:19]
  wire  top_io_out_ar_valid; // @[SimTop.scala 23:19]
  wire [31:0] top_io_out_ar_bits_addr; // @[SimTop.scala 23:19]
  wire  top_io_out_r_ready; // @[SimTop.scala 23:19]
  wire  top_io_out_r_valid; // @[SimTop.scala 23:19]
  wire [63:0] top_io_out_r_bits_data; // @[SimTop.scala 23:19]
  wire  top_io_out_r_bits_last; // @[SimTop.scala 23:19]
  wire  top_io_imem_inst_valid; // @[SimTop.scala 23:19]
  wire  top_io_imem_inst_ready; // @[SimTop.scala 23:19]
  wire [31:0] top_io_imem_inst_addr; // @[SimTop.scala 23:19]
  wire [127:0] top_io_imem_inst_read; // @[SimTop.scala 23:19]
  wire  top_io_dmem_data_valid; // @[SimTop.scala 23:19]
  wire  top_io_dmem_data_ready; // @[SimTop.scala 23:19]
  wire  top_io_dmem_data_req; // @[SimTop.scala 23:19]
  wire [31:0] top_io_dmem_data_addr; // @[SimTop.scala 23:19]
  wire [7:0] top_io_dmem_data_strb; // @[SimTop.scala 23:19]
  wire [127:0] top_io_dmem_data_read; // @[SimTop.scala 23:19]
  wire [127:0] top_io_dmem_data_write; // @[SimTop.scala 23:19]
  Core core ( // @[SimTop.scala 18:20]
    .clock(core_clock),
    .reset(core_reset),
    .io_imem_inst_valid(core_io_imem_inst_valid),
    .io_imem_inst_ready(core_io_imem_inst_ready),
    .io_imem_inst_addr(core_io_imem_inst_addr),
    .io_imem_inst_read(core_io_imem_inst_read),
    .io_dmem_data_valid(core_io_dmem_data_valid),
    .io_dmem_data_ready(core_io_dmem_data_ready),
    .io_dmem_data_req(core_io_dmem_data_req),
    .io_dmem_data_addr(core_io_dmem_data_addr),
    .io_dmem_data_size(core_io_dmem_data_size),
    .io_dmem_data_strb(core_io_dmem_data_strb),
    .io_dmem_data_read(core_io_dmem_data_read),
    .io_dmem_data_write(core_io_dmem_data_write)
  );
  ICache icache ( // @[SimTop.scala 19:22]
    .clock(icache_clock),
    .reset(icache_reset),
    .io_imem_inst_valid(icache_io_imem_inst_valid),
    .io_imem_inst_ready(icache_io_imem_inst_ready),
    .io_imem_inst_addr(icache_io_imem_inst_addr),
    .io_imem_inst_read(icache_io_imem_inst_read),
    .io_out_inst_valid(icache_io_out_inst_valid),
    .io_out_inst_ready(icache_io_out_inst_ready),
    .io_out_inst_addr(icache_io_out_inst_addr),
    .io_out_inst_read(icache_io_out_inst_read)
  );
  DCache dcache ( // @[SimTop.scala 20:22]
    .clock(dcache_clock),
    .reset(dcache_reset),
    .io_dmem_data_valid(dcache_io_dmem_data_valid),
    .io_dmem_data_ready(dcache_io_dmem_data_ready),
    .io_dmem_data_req(dcache_io_dmem_data_req),
    .io_dmem_data_addr(dcache_io_dmem_data_addr),
    .io_dmem_data_size(dcache_io_dmem_data_size),
    .io_dmem_data_strb(dcache_io_dmem_data_strb),
    .io_dmem_data_read(dcache_io_dmem_data_read),
    .io_dmem_data_write(dcache_io_dmem_data_write),
    .io_out_data_valid(dcache_io_out_data_valid),
    .io_out_data_ready(dcache_io_out_data_ready),
    .io_out_data_req(dcache_io_out_data_req),
    .io_out_data_addr(dcache_io_out_data_addr),
    .io_out_data_strb(dcache_io_out_data_strb),
    .io_out_data_read(dcache_io_out_data_read),
    .io_out_data_write(dcache_io_out_data_write)
  );
  AxiLite2Axi top ( // @[SimTop.scala 23:19]
    .clock(top_clock),
    .reset(top_reset),
    .io_out_aw_ready(top_io_out_aw_ready),
    .io_out_aw_valid(top_io_out_aw_valid),
    .io_out_aw_bits_addr(top_io_out_aw_bits_addr),
    .io_out_w_ready(top_io_out_w_ready),
    .io_out_w_valid(top_io_out_w_valid),
    .io_out_w_bits_data(top_io_out_w_bits_data),
    .io_out_w_bits_strb(top_io_out_w_bits_strb),
    .io_out_w_bits_last(top_io_out_w_bits_last),
    .io_out_b_ready(top_io_out_b_ready),
    .io_out_b_valid(top_io_out_b_valid),
    .io_out_ar_ready(top_io_out_ar_ready),
    .io_out_ar_valid(top_io_out_ar_valid),
    .io_out_ar_bits_addr(top_io_out_ar_bits_addr),
    .io_out_r_ready(top_io_out_r_ready),
    .io_out_r_valid(top_io_out_r_valid),
    .io_out_r_bits_data(top_io_out_r_bits_data),
    .io_out_r_bits_last(top_io_out_r_bits_last),
    .io_imem_inst_valid(top_io_imem_inst_valid),
    .io_imem_inst_ready(top_io_imem_inst_ready),
    .io_imem_inst_addr(top_io_imem_inst_addr),
    .io_imem_inst_read(top_io_imem_inst_read),
    .io_dmem_data_valid(top_io_dmem_data_valid),
    .io_dmem_data_ready(top_io_dmem_data_ready),
    .io_dmem_data_req(top_io_dmem_data_req),
    .io_dmem_data_addr(top_io_dmem_data_addr),
    .io_dmem_data_strb(top_io_dmem_data_strb),
    .io_dmem_data_read(top_io_dmem_data_read),
    .io_dmem_data_write(top_io_dmem_data_write)
  );
  assign io_uart_out_valid = 1'h0; // @[SimTop.scala 41:21]
  assign io_uart_out_ch = 8'h0; // @[SimTop.scala 42:18]
  assign io_uart_in_valid = 1'h0; // @[SimTop.scala 43:20]
  assign io_memAXI_0_aw_valid = top_io_out_aw_valid; // @[SimTop.scala 32:18]
  assign io_memAXI_0_aw_bits_addr = top_io_out_aw_bits_addr; // @[SimTop.scala 32:18]
  assign io_memAXI_0_aw_bits_prot = 3'h0; // @[SimTop.scala 32:18]
  assign io_memAXI_0_aw_bits_id = 4'h0; // @[SimTop.scala 32:18]
  assign io_memAXI_0_aw_bits_user = 1'h0; // @[SimTop.scala 32:18]
  assign io_memAXI_0_aw_bits_len = 8'h0; // @[SimTop.scala 32:18]
  assign io_memAXI_0_aw_bits_size = 3'h3; // @[SimTop.scala 32:18]
  assign io_memAXI_0_aw_bits_burst = 2'h1; // @[SimTop.scala 32:18]
  assign io_memAXI_0_aw_bits_lock = 1'h0; // @[SimTop.scala 32:18]
  assign io_memAXI_0_aw_bits_cache = 4'h2; // @[SimTop.scala 32:18]
  assign io_memAXI_0_aw_bits_qos = 4'h0; // @[SimTop.scala 32:18]
  assign io_memAXI_0_w_valid = top_io_out_w_valid; // @[SimTop.scala 33:18]
  assign io_memAXI_0_w_bits_data[0] = top_io_out_w_bits_data; // @[SimTop.scala 33:18]
  assign io_memAXI_0_w_bits_strb = top_io_out_w_bits_strb; // @[SimTop.scala 33:18]
  assign io_memAXI_0_w_bits_last = 1'h1; // @[SimTop.scala 33:18]
  assign io_memAXI_0_b_ready = 1'h1; // @[SimTop.scala 34:18]
  assign io_memAXI_0_ar_valid = top_io_out_ar_valid; // @[SimTop.scala 35:18]
  assign io_memAXI_0_ar_bits_addr = top_io_out_ar_bits_addr; // @[SimTop.scala 35:18]
  assign io_memAXI_0_ar_bits_prot = 3'h0; // @[SimTop.scala 35:18]
  assign io_memAXI_0_ar_bits_id = 4'h0; // @[SimTop.scala 35:18]
  assign io_memAXI_0_ar_bits_user = 1'h0; // @[SimTop.scala 35:18]
  assign io_memAXI_0_ar_bits_len = 8'h1; // @[SimTop.scala 35:18]
  assign io_memAXI_0_ar_bits_size = 3'h3; // @[SimTop.scala 35:18]
  assign io_memAXI_0_ar_bits_burst = 2'h1; // @[SimTop.scala 35:18]
  assign io_memAXI_0_ar_bits_lock = 1'h0; // @[SimTop.scala 35:18]
  assign io_memAXI_0_ar_bits_cache = 4'h2; // @[SimTop.scala 35:18]
  assign io_memAXI_0_ar_bits_qos = 4'h0; // @[SimTop.scala 35:18]
  assign io_memAXI_0_r_ready = 1'h1; // @[SimTop.scala 36:18]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_imem_inst_ready = icache_io_imem_inst_ready; // @[SimTop.scala 27:17]
  assign core_io_imem_inst_read = icache_io_imem_inst_read; // @[SimTop.scala 27:17]
  assign core_io_dmem_data_ready = dcache_io_dmem_data_ready; // @[SimTop.scala 29:17]
  assign core_io_dmem_data_read = dcache_io_dmem_data_read; // @[SimTop.scala 29:17]
  assign icache_clock = clock;
  assign icache_reset = reset;
  assign icache_io_imem_inst_valid = core_io_imem_inst_valid; // @[SimTop.scala 27:17]
  assign icache_io_imem_inst_addr = core_io_imem_inst_addr; // @[SimTop.scala 27:17]
  assign icache_io_out_inst_ready = top_io_imem_inst_ready; // @[SimTop.scala 28:17]
  assign icache_io_out_inst_read = top_io_imem_inst_read; // @[SimTop.scala 28:17]
  assign dcache_clock = clock;
  assign dcache_reset = reset;
  assign dcache_io_dmem_data_valid = core_io_dmem_data_valid; // @[SimTop.scala 29:17]
  assign dcache_io_dmem_data_req = core_io_dmem_data_req; // @[SimTop.scala 29:17]
  assign dcache_io_dmem_data_addr = core_io_dmem_data_addr; // @[SimTop.scala 29:17]
  assign dcache_io_dmem_data_size = core_io_dmem_data_size; // @[SimTop.scala 29:17]
  assign dcache_io_dmem_data_strb = core_io_dmem_data_strb; // @[SimTop.scala 29:17]
  assign dcache_io_dmem_data_write = core_io_dmem_data_write; // @[SimTop.scala 29:17]
  assign dcache_io_out_data_ready = top_io_dmem_data_ready; // @[SimTop.scala 30:17]
  assign dcache_io_out_data_read = top_io_dmem_data_read; // @[SimTop.scala 30:17]
  assign top_clock = clock;
  assign top_reset = reset;
  assign top_io_out_aw_ready = io_memAXI_0_aw_ready; // @[SimTop.scala 32:18]
  assign top_io_out_w_ready = io_memAXI_0_w_ready; // @[SimTop.scala 33:18]
  assign top_io_out_b_valid = io_memAXI_0_b_valid; // @[SimTop.scala 34:18]
  assign top_io_out_ar_ready = io_memAXI_0_ar_ready; // @[SimTop.scala 35:18]
  assign top_io_out_r_valid = io_memAXI_0_r_valid; // @[SimTop.scala 36:18]
  assign top_io_out_r_bits_data = io_memAXI_0_r_bits_data[0]; // @[SimTop.scala 36:18]
  assign top_io_out_r_bits_last = io_memAXI_0_r_bits_last; // @[SimTop.scala 36:18]
  assign top_io_imem_inst_valid = icache_io_out_inst_valid; // @[SimTop.scala 28:17]
  assign top_io_imem_inst_addr = icache_io_out_inst_addr; // @[SimTop.scala 28:17]
  assign top_io_dmem_data_valid = dcache_io_out_data_valid; // @[SimTop.scala 30:17]
  assign top_io_dmem_data_req = dcache_io_out_data_req; // @[SimTop.scala 30:17]
  assign top_io_dmem_data_addr = dcache_io_out_data_addr; // @[SimTop.scala 30:17]
  assign top_io_dmem_data_strb = dcache_io_out_data_strb; // @[SimTop.scala 30:17]
  assign top_io_dmem_data_write = dcache_io_out_data_write; // @[SimTop.scala 30:17]
endmodule
